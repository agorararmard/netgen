* NGSPICE file created from xtea.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 D Q RESET_B CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

.subckt xtea all_done clock data_in1[0] data_in1[10] data_in1[11] data_in1[12] data_in1[13]
+ data_in1[14] data_in1[15] data_in1[16] data_in1[17] data_in1[18] data_in1[19] data_in1[1]
+ data_in1[20] data_in1[21] data_in1[22] data_in1[23] data_in1[24] data_in1[25] data_in1[26]
+ data_in1[27] data_in1[28] data_in1[29] data_in1[2] data_in1[30] data_in1[31] data_in1[3]
+ data_in1[4] data_in1[5] data_in1[6] data_in1[7] data_in1[8] data_in1[9] data_in2[0]
+ data_in2[10] data_in2[11] data_in2[12] data_in2[13] data_in2[14] data_in2[15] data_in2[16]
+ data_in2[17] data_in2[18] data_in2[19] data_in2[1] data_in2[20] data_in2[21] data_in2[22]
+ data_in2[23] data_in2[24] data_in2[25] data_in2[26] data_in2[27] data_in2[28] data_in2[29]
+ data_in2[2] data_in2[30] data_in2[31] data_in2[3] data_in2[4] data_in2[5] data_in2[6]
+ data_in2[7] data_in2[8] data_in2[9] data_out1[0] data_out1[10] data_out1[11] data_out1[12]
+ data_out1[13] data_out1[14] data_out1[15] data_out1[16] data_out1[17] data_out1[18]
+ data_out1[19] data_out1[1] data_out1[20] data_out1[21] data_out1[22] data_out1[23]
+ data_out1[24] data_out1[25] data_out1[26] data_out1[27] data_out1[28] data_out1[29]
+ data_out1[2] data_out1[30] data_out1[31] data_out1[3] data_out1[4] data_out1[5]
+ data_out1[6] data_out1[7] data_out1[8] data_out1[9] data_out2[0] data_out2[10] data_out2[11]
+ data_out2[12] data_out2[13] data_out2[14] data_out2[15] data_out2[16] data_out2[17]
+ data_out2[18] data_out2[19] data_out2[1] data_out2[20] data_out2[21] data_out2[22]
+ data_out2[23] data_out2[24] data_out2[25] data_out2[26] data_out2[27] data_out2[28]
+ data_out2[29] data_out2[2] data_out2[30] data_out2[31] data_out2[3] data_out2[4]
+ data_out2[5] data_out2[6] data_out2[7] data_out2[8] data_out2[9] key_in[0] key_in[100]
+ key_in[101] key_in[102] key_in[103] key_in[104] key_in[105] key_in[106] key_in[107]
+ key_in[108] key_in[109] key_in[10] key_in[110] key_in[111] key_in[112] key_in[113]
+ key_in[114] key_in[115] key_in[116] key_in[117] key_in[118] key_in[119] key_in[11]
+ key_in[120] key_in[121] key_in[122] key_in[123] key_in[124] key_in[125] key_in[126]
+ key_in[127] key_in[12] key_in[13] key_in[14] key_in[15] key_in[16] key_in[17] key_in[18]
+ key_in[19] key_in[1] key_in[20] key_in[21] key_in[22] key_in[23] key_in[24] key_in[25]
+ key_in[26] key_in[27] key_in[28] key_in[29] key_in[2] key_in[30] key_in[31] key_in[32]
+ key_in[33] key_in[34] key_in[35] key_in[36] key_in[37] key_in[38] key_in[39] key_in[3]
+ key_in[40] key_in[41] key_in[42] key_in[43] key_in[44] key_in[45] key_in[46] key_in[47]
+ key_in[48] key_in[49] key_in[4] key_in[50] key_in[51] key_in[52] key_in[53] key_in[54]
+ key_in[55] key_in[56] key_in[57] key_in[58] key_in[59] key_in[5] key_in[60] key_in[61]
+ key_in[62] key_in[63] key_in[64] key_in[65] key_in[66] key_in[67] key_in[68] key_in[69]
+ key_in[6] key_in[70] key_in[71] key_in[72] key_in[73] key_in[74] key_in[75] key_in[76]
+ key_in[77] key_in[78] key_in[79] key_in[7] key_in[80] key_in[81] key_in[82] key_in[83]
+ key_in[84] key_in[85] key_in[86] key_in[87] key_in[88] key_in[89] key_in[8] key_in[90]
+ key_in[91] key_in[92] key_in[93] key_in[94] key_in[95] key_in[96] key_in[97] key_in[98]
+ key_in[99] key_in[9] mode reset VPWR VGND
XFILLER_79_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_918 VGND VPWR sky130_fd_sc_hd__decap_12
X_3155_ _3155_/A _3155_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4935__A _4642_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_277 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_586 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_512 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_737 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_372 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_748 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_383 VGND VPWR sky130_fd_sc_hd__fill_2
X_3086_ _2943_/A _4043_/C _3875_/A _3253_/A _3087_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4654__B _4586_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_545 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_770 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_589 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_280 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_965 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_628 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_818 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4670__A _4527_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_166 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5196__A2 _4574_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3988_ _3903_/X _3964_/X _3988_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_497 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_801 VGND VPWR sky130_fd_sc_hd__decap_12
X_2939_ _2931_/Y _2938_/X _2931_/Y _2938_/X _2939_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_834 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3717__C _3716_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_4609_ _4646_/B _4609_/B _4609_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_116_260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_720 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_794 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3201__A1_N _3188_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_111 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3733__B _3727_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_466 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_797 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_959 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3534__B1_N _3507_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5503__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_661 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3846__A1_N _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_748 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4564__B _4561_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2890__B1 _5261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_483 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_239 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__C1 _4918_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4580__A _5256_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_678 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_464 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5187__A2 key_in[96] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2812__B _2698_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_672 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3196__A _3124_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_683 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_311 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_867 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_837 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3924__A _3895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5561__D _4559_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_572 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_937 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3362__C _3362_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_637 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5111__A2 _5108_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_531 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3122__A1 _4638_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_851 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3122__B2 _3121_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_545 VGND VPWR sky130_fd_sc_hd__decap_8
X_4960_ _4947_/X _4950_/X _4960_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_18_984 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3425__A2 _3421_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_781 VGND VPWR sky130_fd_sc_hd__decap_12
X_3911_ _3861_/X _3891_/X _3864_/Y _3912_/C VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_17_494 VGND VPWR sky130_fd_sc_hd__fill_2
X_4891_ _4891_/A _4889_/Y _4890_/X _4891_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4490__A _4269_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3842_ _3721_/Y _3841_/X _3842_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_60_784 VGND VPWR sky130_fd_sc_hd__decap_3
X_3773_ _3769_/Y _3771_/X _3819_/A _3773_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__2722__B _2722_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2936__A1 _4637_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_823 VGND VPWR sky130_fd_sc_hd__fill_1
X_5512_ _5220_/X _3588_/A _4348_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2936__B2 _2935_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2724_ _2723_/A _2723_/B _2776_/A _2728_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_157_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_693 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_181 VGND VPWR sky130_fd_sc_hd__decap_3
X_5443_ _5443_/D _5443_/Q _4430_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4689__A1 _5356_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4689__B2 _4688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_837 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3834__A _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5374_ _5374_/D data_out1[4] _4512_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4649__B _4523_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_369 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5526__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_4325_ _4324_/A _4325_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5471__D _5089_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3645__A2_N _3644_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_594 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_4256_ _4256_/A _4658_/X _4256_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_102_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_3207_ _3143_/C _3166_/B _3207_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4665__A _4664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_350 VGND VPWR sky130_fd_sc_hd__decap_12
X_4187_ _4073_/X _4187_/B _4187_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_68_884 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4861__A1 _5548_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_832 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_383 VGND VPWR sky130_fd_sc_hd__decap_12
X_3138_ _3135_/X _3137_/Y _3138_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_82_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_68 VGND VPWR sky130_fd_sc_hd__fill_2
X_3069_ _3069_/A _3068_/Y _3071_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_24_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_515 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4613__B2 _4610_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_420 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_239 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_453 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2913__A _2913_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_615 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3728__B _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_125 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_536 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_152 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_54 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_686 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3744__A _3743_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4559__B _4557_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_742 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_69 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5381__D _4761_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4575__A _4518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_737 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_128 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2863__B1 _2861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_62 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_84 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_898 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4604__A1 _5443_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_921 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_537 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_559 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4080__A2 _4055_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_913 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_998 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_250 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_83 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_283 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3638__B _3638_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_94 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5556__D _4553_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5549__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3591__B2 _3590_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5547__RESET_B _4306_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3654__A _3615_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3738__A1_N _3720_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5119__A2_N _5118_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_615 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_892 VGND VPWR sky130_fd_sc_hd__decap_4
X_4110_ _4109_/X _4152_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_78_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_957 VGND VPWR sky130_fd_sc_hd__decap_12
X_5090_ _5472_/Q _5090_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_158 VGND VPWR sky130_fd_sc_hd__fill_1
X_4041_ _3974_/A _4041_/B _4041_/C _4041_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4485__A _4483_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_810 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_117 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3820__C _3774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_534 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2717__B _2717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_813 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_161 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_172 VGND VPWR sky130_fd_sc_hd__fill_1
X_4943_ _4943_/A _4943_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4932__B _4922_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3829__A _3829_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2733__A _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_773 VGND VPWR sky130_fd_sc_hd__fill_1
X_4874_ _4874_/A _4873_/Y _4874_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_21_935 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_929 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_434 VGND VPWR sky130_fd_sc_hd__decap_4
X_3825_ _3815_/Y _3824_/Y _3815_/Y _3824_/Y _3825_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5466__D _5022_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3756_ _2796_/X _3755_/X _2796_/X _3755_/X _3756_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3031__B1 _2714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_642 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_333 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2947__A1_N _2939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_867 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5244__A1_N _5227_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2707_ _2707_/A key_in[71] _2707_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_601 VGND VPWR sky130_fd_sc_hd__fill_1
X_3687_ _3685_/X _3686_/Y _3687_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_837 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3564__A _3564_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_528 VGND VPWR sky130_fd_sc_hd__decap_3
X_5426_ _5426_/D data_out2[24] _4451_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3283__B _3282_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5357_ _5323_/X _5347_/Y _5357_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_188 VGND VPWR sky130_fd_sc_hd__decap_12
X_4308_ _4305_/A _4308_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_391 VGND VPWR sky130_fd_sc_hd__fill_2
X_5288_ _5288_/A _2799_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_88_979 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_169 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4395__A _4390_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4239_ _3397_/Y _3556_/Y _3397_/Y _3556_/Y _4239_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_266 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2908__A _2832_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_489 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3637__A2 _5520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_990 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_45 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2845__B1 _2844_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_802 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_684 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_44 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4598__B1 _4597_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4842__B _4842_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4062__A2 _4058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_902 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3739__A _5292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_913 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_423 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3458__B _3459_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_255 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_979 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5376__D _4751_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3537__A2_N _3536_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_489 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_97 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_46 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_611 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_358 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3094__A1_N _3176_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3876__A2 _3875_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_968 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_456 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3921__B _3921_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3089__B1 _3088_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2836__B1 _2794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_813 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_150 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_684 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3649__A _3626_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_378 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_929 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5371__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_3610_ _3583_/C _3593_/X _3595_/X _3610_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
X_4590_ _4590_/A _4590_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_128_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_804 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4761__B1 data_out1[11] VGND VPWR sky130_fd_sc_hd__diode_2
X_3541_ _3489_/A _3513_/A _3541_/C _3541_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_156_984 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_163 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5381__RESET_B _4503_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_196 VGND VPWR sky130_fd_sc_hd__decap_8
X_3472_ _3501_/A key_in[92] _3472_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5305__A2 _5300_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4199__B _4198_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5211_ _5211_/A _5210_/X _5211_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_306 VGND VPWR sky130_fd_sc_hd__fill_1
X_5142_ _4857_/A _5139_/X _5141_/Y _5128_/A _4815_/A _5142_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_111_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_754 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4927__B _4917_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_242 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3831__B _3829_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_916 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2728__A _2728_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5073_ _5071_/Y _5072_/X _4803_/Y _5073_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_56_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_629 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4816__A1 _4802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4646__C _5446_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5104__A _5104_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4816__B2 _4815_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4024_ _3974_/A _4027_/B _4024_/C _4024_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_84_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_971 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4943__A _4943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_684 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_345 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4662__B _4586_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_654 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_4926_ _4925_/A _4924_/X _4925_/X _4928_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3252__B1 _5497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4857_ _4857_/A _4855_/X _4856_/Y _4857_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_21_765 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5469__RESET_B _4399_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_759 VGND VPWR sky130_fd_sc_hd__decap_4
X_3808_ _3791_/Y _3806_/X _3808_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3004__B1 _3002_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_951 VGND VPWR sky130_fd_sc_hd__decap_8
X_4788_ _3178_/A _4788_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_153_409 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_130 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4752__B1 data_out1[7] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3555__B2 _3554_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_601 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2910__B _2908_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3739_ _5292_/X _3738_/X _3739_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_109_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_483 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_623 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_27 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_38 VGND VPWR sky130_fd_sc_hd__fill_2
X_5409_ _4690_/X data_out2[7] _4471_/X _5402_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3307__B2 _3306_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4820__A2_N _4819_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_614 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_754 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4837__B _4837_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3741__B _3713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_275 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4807__A1 _4798_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4807__B2 _4806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5014__A _4559_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3460__C _3460_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_843 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_331 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2818__B1 _4750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_876 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_64 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_643 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4572__B _4561_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5394__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3469__A _3469_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_367 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4035__A2 _4011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5232__B2 _5201_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_743 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_417 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_707 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_951 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_235 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3546__A1 data_in2[30] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_257 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3916__B _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_910 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_268 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4743__B1 data_out1[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_931 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_997 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3849__A2 _3824_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3932__A _4720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1016 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_618 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3651__B _3649_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_938 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_640 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4763__A _2737_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_846 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_507 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3379__A _5472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_985 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_687 VGND VPWR sky130_fd_sc_hd__fill_2
X_2972_ _4637_/X _2968_/X _2969_/X _2970_/X _2971_/X _2972_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_43_890 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4711_ _3073_/C _4699_/X data_out2[17] _4701_/X _5419_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3098__B _3099_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5562__RESET_B _4288_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4642_ _4642_/A _4642_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3826__B _3825_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_729 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3537__B2 _3536_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4573_ _4573_/A _4561_/B _4573_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_129_995 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_3524_ _3396_/X _3523_/X _3396_/X _3523_/X _3526_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_791 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3545__C _3545_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_144 VGND VPWR sky130_fd_sc_hd__decap_12
X_3455_ _4731_/X _3455_/B _3488_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_103_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4938__A _4938_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3842__A _3721_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4657__B _4522_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3386_ _4728_/X _3385_/B _3385_/X _3388_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3242__B1_N _3241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3561__B _3561_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_5125_ _5125_/A _5124_/X _5125_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_873 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_117 VGND VPWR sky130_fd_sc_hd__decap_4
X_5056_ _5056_/A _5056_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_66_960 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4265__A2 _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_982 VGND VPWR sky130_fd_sc_hd__decap_3
X_4007_ _3959_/X _4007_/B _4007_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4673__A _4672_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3473__B1 _3408_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_846 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_857 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5214__B2 _5213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_676 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3289__A _3249_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_501 VGND VPWR sky130_fd_sc_hd__decap_6
X_4909_ _4873_/A _4908_/X _4909_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3776__B2 _3775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4973__B1 _5462_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_562 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2921__A _2850_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_205 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_623 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5009__A _5008_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_965 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_902 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4848__A _4848_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_486 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3752__A _3636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_979 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4567__B _4557_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3471__B key_in[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_466 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_949 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_919 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_802 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_109 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_418 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_813 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4583__A _4582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_492 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2815__B _2814_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3199__A _3199_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_698 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_340 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_871 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3927__A _3835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2831__A _4907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2990__A2 _2989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4716__B1 data_out2[19] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5564__D _4563_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_45 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_559 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4192__B2 _4191_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_475 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2742__A2 _2739_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4758__A _4701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3662__A _5516_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_3240_ _3249_/B _3239_/X _3249_/B _3239_/X _3280_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_136 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4908__D _5552_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_713 VGND VPWR sky130_fd_sc_hd__fill_2
X_3171_ data_in2[19] _2956_/X _3143_/X _3170_/Y _3171_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_94_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4247__A2 _4246_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_204 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4493__A _4492_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_470 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_259 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_602 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5101__B _5091_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_646 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3758__B2 _3757_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2955_ data_in2[13] _2731_/X _2929_/X _2954_/Y _5524_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4940__B _4938_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_860 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3837__A _4533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3306__A2_N _3305_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2741__A _2741_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_370 VGND VPWR sky130_fd_sc_hd__decap_12
X_2886_ _5523_/Q _2918_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_163_504 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3556__B _3555_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4625_ _3148_/A _3293_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_129_770 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5474__D _5127_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4556_ _4546_/A _4557_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_442 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_913 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_773 VGND VPWR sky130_fd_sc_hd__decap_12
X_3507_ _3505_/X _3507_/B _3507_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_998 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_208 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4668__A _4667_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_315 VGND VPWR sky130_fd_sc_hd__decap_3
X_4487_ _4483_/X _4487_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3572__A _5516_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3181__B1_N _3236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_114 VGND VPWR sky130_fd_sc_hd__decap_8
X_3438_ _3465_/A _3464_/A _3438_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_103_136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_979 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3291__B key_in[55] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_489 VGND VPWR sky130_fd_sc_hd__decap_4
X_3369_ _3233_/A _3368_/A _4778_/X _3368_/Y _3369_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_5108_ _5087_/A _5098_/A _5108_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_245 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4238__A2 _4228_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_418 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_278 VGND VPWR sky130_fd_sc_hd__fill_1
X_5039_ _5037_/X _5038_/X _5039_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_598 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2916__A _2998_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3446__B1 _3408_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_492 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_67 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_985 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5484__RESET_B _4381_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5011__B _5007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_495 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5413__RESET_B _4466_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_309 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_292 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4946__B1 _4553_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4850__B _4849_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_98 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5432__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_567 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_887 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3466__B _3466_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2972__A2 _2968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_514 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5384__D _4766_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_559 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_75 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2724__A2 _2723_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4578__A _4578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4083__A2_N _4082_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3482__A _3463_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_753 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_370 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_908 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_513 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2826__A _2861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_440 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5559__D _5559_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_473 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_646 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_820 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__A _3634_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_831 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_189 VGND VPWR sky130_fd_sc_hd__fill_2
X_2740_ _2740_/A _2741_/A VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4036__A2_N _4035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3376__B key_in[89] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_396 VGND VPWR sky130_fd_sc_hd__fill_1
X_4410_ _4411_/A _4410_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5390_ _4777_/X data_out1[20] _4493_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_126_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_913 VGND VPWR sky130_fd_sc_hd__decap_3
X_4341_ _4341_/A _4341_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2715__A2 _2714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_261 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4488__A _4483_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_635 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3392__A _5223_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_294 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_231 VGND VPWR sky130_fd_sc_hd__fill_2
X_4272_ _4271_/A _4272_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_979 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1009 VGND VPWR sky130_fd_sc_hd__decap_8
X_3223_ _3291_/A key_in[117] _3222_/X _3223_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_98_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_521 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_117 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_128 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_841 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_3154_ _3197_/B _3153_/Y _3197_/B _3153_/Y _3154_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4935__B _4934_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_524 VGND VPWR sky130_fd_sc_hd__fill_2
X_3085_ _3085_/A _3253_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3230__A2_N _3229_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_535 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3428__B1 _3385_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5112__A _5113_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4654__C _4519_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_248 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5469__D _5063_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_782 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4951__A _4951_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5455__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_977 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4670__B _4616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3987_ _3154_/X _3986_/X _3154_/X _3986_/X _3987_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_843 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_15_0_clock clkbuf_3_7_0_clock/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_329 VGND VPWR sky130_fd_sc_hd__decap_6
X_2938_ _4943_/A _2936_/X _2937_/X _2938_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_164_813 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_312 VGND VPWR sky130_fd_sc_hd__fill_2
X_2869_ _2870_/A _2870_/B _2871_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4176__A1_N _3452_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_4608_ _4646_/A _4605_/B _4607_/Y _5444_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_163_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_762 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4398__A _4402_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4539_ _5197_/A _4541_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_743 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_957 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_968 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_294 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3733__C _3731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_445 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_89 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_478 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_532 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_204 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_673 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_790 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2890__A1 _5292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2890__B2 _2889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5379__D _4755_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_86 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_590 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__B1 _4531_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_476 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3477__A _3475_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_30 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_41 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_651 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2812__C _2842_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3196__B _3196_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_537 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4147__A1 _3395_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_333 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3924__B _3920_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_399 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4101__A _4100_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_46 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_949 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_521 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_148 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3122__A2 _3118_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_321 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_941 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5478__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_343 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4083__B1 _4075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3910_ _3860_/X _3888_/X _3910_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4890_ _4886_/X _4888_/X _4890_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_32_421 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_281 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5349__A2_N _5348_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3841_ _3636_/Y _5529_/Q _2847_/A _3133_/A _3841_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_33_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3387__A _3388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_3 VGND VPWR sky130_fd_sc_hd__decap_8
X_3772_ _3769_/Y _3771_/X _3819_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_121_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2936__A2 _2932_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2723_ _2723_/A _2723_/B _2776_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_5511_ _5196_/X _3573_/A _4349_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_9_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_857 VGND VPWR sky130_fd_sc_hd__decap_4
X_5442_ _4599_/Y _4600_/A _4431_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_118_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4689__A2 _4687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_378 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3834__B _3832_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5373_ _5373_/D data_out1[3] _4513_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_126_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_4324_ _4324_/A _4324_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_231 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_776 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_415 VGND VPWR sky130_fd_sc_hd__decap_8
X_4255_ _4631_/Y _4264_/B _4255_/C _4254_/X _4255_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3609__B1_N _3608_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_275 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1003 VGND VPWR sky130_fd_sc_hd__fill_2
X_3206_ _3135_/X _3209_/B _3206_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4186_ _4170_/X _4176_/Y _4187_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_971 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2865__B1_N _2864_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4861__A2 _4849_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3137_ _3074_/A _3096_/X _3136_/X _3137_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_95_693 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_237 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_855 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_3068_ _3021_/A _3064_/Y _3066_/Y _3067_/Y _3068_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_55_579 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_922 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_782 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_955 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_605 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_465 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2913__B _2912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3728__C _3706_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_695 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_345 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5326__B1 _5199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_815 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5017__A _5017_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_551 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_787 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4856__A _4853_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_841 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4575__B _4524_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_885 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_671 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_384 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2863__A1 _4637_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2863__B2 _2862_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_708 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_64 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4065__B1 _4037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4604__A2 _4601_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_229 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4591__A _4590_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_51 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_988 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_487 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_796 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_95 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3000__A _2898_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3935__A _5528_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_868 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_879 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_367 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3654__B _3570_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5572__D _4572_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_697 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_174 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_197 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_562 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_627 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_947 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_892 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_969 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3670__A _3658_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5516__RESET_B _4343_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_4040_ _4039_/A _4038_/X _4041_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_1_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5273__A2_N _5272_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4969__B1_N _4968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_4942_ _4546_/A _4942_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3803__B1 _3794_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_292 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3829__B _3806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2733__B _2698_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4873_ _4873_/A _4872_/X _4873_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_32_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_571 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4006__A _3961_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3824_ _3823_/X _3824_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_159_993 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_301 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_824 VGND VPWR sky130_fd_sc_hd__decap_12
X_3755_ _3753_/X _3754_/X _3755_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__3031__A1 _2714_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3031__B2 _3233_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5308__B1 _5270_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2706_ _5236_/A key_in[7] _2706_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_805 VGND VPWR sky130_fd_sc_hd__fill_1
X_3686_ _3661_/X _3667_/X _3663_/X _3686_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_145_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_624 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3564__B _3564_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_849 VGND VPWR sky130_fd_sc_hd__decap_12
X_5425_ _5425_/D data_out2[23] _4452_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5482__D _3632_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_5356_ _5252_/A _2698_/B _5356_/C _5356_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_0_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_18 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_273 VGND VPWR sky130_fd_sc_hd__decap_8
X_4307_ _4305_/A _4307_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_947 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4676__A _4700_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5287_ _5287_/A _5290_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_59_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_234 VGND VPWR sky130_fd_sc_hd__fill_2
X_4238_ _3523_/X _4228_/X _4236_/B _4246_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_101_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_479 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2908__B _2864_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_278 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_693 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_129 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2845__A1 _2842_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4169_ _4151_/X _4170_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_74_17 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_321 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_505 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_527 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4598__A1 _5441_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_538 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2924__A _2878_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_869 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5300__A _5300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3739__B _3738_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_240 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_223 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_947 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_593 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_407 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_109 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_406 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_417 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3755__A _3753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_602 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_304 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3691__A2_N _3690_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5392__D _5392_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_690 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4586__A _4524_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_199 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3490__A _3489_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3089__A1 _2889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_479 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2836__A1 _2761_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_365 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_538 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2834__A _2762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_752 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_357 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3649__B _3631_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5567__D _4566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5516__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_295 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_788 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4210__B1 _4208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3665__A _3661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_940 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4761__A1 _3804_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3540_ _3540_/A _3540_/B _3540_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_143_602 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4761__B2 _4758_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_816 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_450 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3659__A2_N _5521_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2772__B1 _2753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_112 VGND VPWR sky130_fd_sc_hd__fill_2
X_3471_ _3501_/A key_in[28] _3471_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_6_483 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5305__A3 _5301_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_657 VGND VPWR sky130_fd_sc_hd__fill_2
X_5210_ _4811_/A _5209_/Y _4811_/A _5209_/Y _5210_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_167 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_413 VGND VPWR sky130_fd_sc_hd__fill_2
X_5141_ _5148_/B _5141_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_510 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4496__A _4492_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_766 VGND VPWR sky130_fd_sc_hd__decap_8
X_5072_ _5072_/A _5072_/B _5072_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_479 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2728__B _2728_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_416 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4816__A2 _4823_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4023_ _4014_/X _4021_/X _4024_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4646__D _4645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5104__B _5103_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4831__B1_N _4830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_505 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2744__A _5332_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_590 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5120__A _5121_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4662__C _4519_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_357 VGND VPWR sky130_fd_sc_hd__decap_8
X_4925_ _4925_/A _4924_/X _4925_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3252__A1 _3110_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5477__D _5477_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3252__B2 _3251_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_908 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_733 VGND VPWR sky130_fd_sc_hd__decap_4
X_4856_ _4853_/X _4854_/X _4856_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3154__A1_N _3197_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3807_ _3791_/Y _3806_/X _3807_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3004__A1 _4637_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3004__B2 _3003_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_276 VGND VPWR sky130_fd_sc_hd__decap_8
X_4787_ _4786_/X _4781_/X data_out1[24] _4782_/X _4787_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_147_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4752__A1 _5229_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_451 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4752__B2 _4746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_816 VGND VPWR sky130_fd_sc_hd__fill_2
X_3738_ _3720_/Y _3737_/X _3720_/Y _3737_/X _3738_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__2910__C _2909_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_996 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_613 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_304 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_687 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_175 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_646 VGND VPWR sky130_fd_sc_hd__decap_12
X_3669_ _3665_/X _3668_/X _3665_/X _3668_/X _3669_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5438__RESET_B _4436_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5408_ _4689_/X data_out2[6] _4472_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_476 VGND VPWR sky130_fd_sc_hd__decap_6
X_5339_ _5299_/A key_in[101] _5303_/A _5339_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4837__C _4541_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_788 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4807__A2 _4813_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5014__B _4997_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_287 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_438 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5103__A2_N _5102_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2818__A1 _5361_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_855 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2818__B2 _3012_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_814 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_674 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_983 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_482 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5539__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_493 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_99 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3737__A1_N _2771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5030__A _5034_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_655 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_143 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3469__B _3468_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_154 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5387__D _4773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_232 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_254 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_930 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3485__A _3431_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4743__A1 _5481_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3546__A2 _3391_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_900 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4743__B2 _4737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_164 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_966 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_420 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_871 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_392 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_906 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_766 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5205__A _4618_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_213 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_747 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_909 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_652 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2946__A1_N _2964_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_814 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_983 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5243__A1_N _5233_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4957__A2_N _4956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_666 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3379__B _3379_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2971_ _2859_/A key_in[110] _2828_/X _2971_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_90_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_699 VGND VPWR sky130_fd_sc_hd__decap_3
X_4710_ _5528_/Q _3073_/C VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4641_ _4640_/X _4631_/Y _5448_/Q _4631_/A _4641_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3395__A _3394_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4572_ _4572_/A _4561_/B _4572_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_613 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_410 VGND VPWR sky130_fd_sc_hd__fill_2
X_3523_ _3368_/Y _3523_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_955 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_443 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5531__RESET_B _4325_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3454_ _3438_/Y _3464_/B _3438_/Y _3464_/B _3455_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_156 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4938__B _4937_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3842__B _3841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_830 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2739__A _5292_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3385_ _4728_/X _3385_/B _3385_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_340 VGND VPWR sky130_fd_sc_hd__fill_2
X_5124_ _5124_/A _5114_/C _5124_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_574 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3536__A2_N _3535_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5055_ _5054_/A _5054_/B _5072_/A _5059_/A VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_69_298 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_758 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4954__A _2973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_4006_ _3961_/Y _4007_/B _4006_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_66_972 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_460 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_825 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3473__A1 _3499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_696 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_324 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_964 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_817 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3289__B _3273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_379 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_828 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_165 VGND VPWR sky130_fd_sc_hd__decap_12
X_4908_ _4874_/A _4872_/X _4908_/C _5552_/Q _4908_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_139_705 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4973__A1 _4870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4973__B2 _4930_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2921__B _2921_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4839_ _5547_/Q _4838_/Y _4839_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_21_596 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_451 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_462 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_229 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2736__B1 _5358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_228 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_605 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_999 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3752__B _3751_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_498 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_968 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5025__A _4975_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_148 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3161__B1 _3183_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_928 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_478 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_585 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_362 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_224 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4864__A _4863_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_65 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_717 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_847 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_869 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_817 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3199__B _3198_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_96 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_330 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_373 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3927__B _3925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_51 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2831__B _2830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_708 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4716__A1 _3143_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4716__B2 _4713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4104__A _4052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_57 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_806 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3943__A _3113_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_251 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_947 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3662__B _3659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_541 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_159 VGND VPWR sky130_fd_sc_hd__decap_8
X_3170_ _3170_/A _3170_/B _3170_/C _3170_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_39_405 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_693 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_555 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_644 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_614 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_997 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_839 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_327 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_658 VGND VPWR sky130_fd_sc_hd__fill_1
X_2954_ _2927_/A _2952_/Y _2953_/X _2954_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4940__C _4949_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2885_ _2885_/A _2927_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_30_382 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_760 VGND VPWR sky130_fd_sc_hd__decap_4
X_4624_ _3077_/A _3148_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_933 VGND VPWR sky130_fd_sc_hd__fill_2
X_4555_ _4555_/A _4541_/B _4555_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4949__A _4949_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3853__A _3840_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_977 VGND VPWR sky130_fd_sc_hd__fill_2
X_3506_ _5128_/A _3474_/X _3477_/X _3507_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_104_605 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_616 VGND VPWR sky130_fd_sc_hd__fill_2
X_4486_ _4483_/X _4486_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_132_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5384__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5490__D _3810_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3437_ _3419_/A _3419_/B _3319_/B _3436_/Y _3464_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_103_148 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_800 VGND VPWR sky130_fd_sc_hd__fill_1
X_3368_ _3368_/A _3368_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3475__A2_N _3474_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_371 VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_clock clkbuf_3_5_0_clock/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_112_682 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_693 VGND VPWR sky130_fd_sc_hd__decap_8
X_5107_ _5104_/A _5103_/X _5124_/A _5113_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4684__A _5516_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3299_ _3297_/X _3298_/Y _3297_/X _3298_/Y _3299_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_58_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_192 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_706 VGND VPWR sky130_fd_sc_hd__fill_2
X_5038_ _5563_/Q _5024_/X _5038_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_899 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_24 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3446__A1 _3499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4643__B1 _4642_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_46 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_143 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_452 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5011__C _5019_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_794 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2932__A _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_658 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4946__B2 _4945_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_833 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_332 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5453__RESET_B _4418_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_708 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_365 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_719 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2972__A3 _2969_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_54 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2709__B1 _2707_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4859__A _4859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_292 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3763__A _3788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_903 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3382__B1 _3414_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_988 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_98 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4578__B _5172_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_284 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3482__B _3482_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3134__B1 _3144_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_765 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_242 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3685__A1 _3589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4594__A _5440_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_728 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2826__B key_in[74] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_611 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4634__B1 _2907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_644 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1000 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_964 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_986 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_772 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_485 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3938__A _3931_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2842__A _2842_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2948__B1 _2888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_310 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_171 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__B _3657_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_182 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_894 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5575__D _4255_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_335 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5362__A1 _5361_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4769__A _4672_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3673__A _3647_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3373__B1 _3371_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4340_ _4340_/A _4341_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_153_571 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_722 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_413 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_582 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_647 VGND VPWR sky130_fd_sc_hd__decap_6
X_4271_ _4271_/A _4271_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_457 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3125__B1 _3124_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_608 VGND VPWR sky130_fd_sc_hd__fill_2
X_3222_ _3044_/X _3222_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_140_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_533 VGND VPWR sky130_fd_sc_hd__decap_12
X_3153_ _3125_/Y _3129_/Y _3124_/Y _3153_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_39_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_706 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3428__A1 _3366_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3084_ _3128_/B _3083_/Y _3128_/B _3083_/Y _3937_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_599 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_227 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5112__B _5111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4654__D _4666_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_290 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4009__A _4003_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_452 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_474 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_625 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_794 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4951__B _4949_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_647 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3848__A _3587_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_433 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2752__A _2752_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4670__C _4661_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3986_ _3984_/X _3985_/X _3984_/X _3985_/X _3986_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_833 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_308 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2939__B1 _2931_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5485__D _3696_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2937_ _4943_/A _2936_/X _2937_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_109_719 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_899 VGND VPWR sky130_fd_sc_hd__fill_2
X_2868_ _2717_/A _3902_/C _5229_/A _3032_/A _2870_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_148_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_858 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_335 VGND VPWR sky130_fd_sc_hd__fill_2
X_4607_ _4609_/B _4607_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4679__A _3588_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2799_ _2799_/A _2799_/B _2799_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3583__A _3615_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_507 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_914 VGND VPWR sky130_fd_sc_hd__fill_1
X_4538_ _4537_/X _5197_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_785 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_936 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_35 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_593 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3733__D _3732_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_809 VGND VPWR sky130_fd_sc_hd__decap_12
X_4469_ _4469_/A _4475_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_917 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_939 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2927__A _2927_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5303__A _5303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_739 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_685 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2890__A2 _2889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_49 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_569 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_43 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_901 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_463 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_608 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_98 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__A1 _4907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_129 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3477__B _3477_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5395__D _5395_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_847 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4147__A2 _4145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4589__A _4589_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3493__A _3519_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_508 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_367 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3924__C _3922_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_880 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_711 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_755 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_809 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_906 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_928 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_544 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3122__A3 _3119_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_330 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5213__A _5212_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_577 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4851__A1_N _5548_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_834 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4083__B2 _4082_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_794 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3668__A _5346_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5375__RESET_B _4510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_433 VGND VPWR sky130_fd_sc_hd__decap_8
X_3840_ _3826_/Y _3833_/Y _3840_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_60_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_606 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_797 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3387__B _3388_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3771_ _3589_/Y _3020_/A _5356_/C _3770_/Y _3771_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_146_803 VGND VPWR sky130_fd_sc_hd__fill_2
X_5510_ _4249_/Y _5510_/Q _4350_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3594__B1 _3583_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2722_ _2722_/A _2722_/B _2723_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__2936__A3 _2933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_184 VGND VPWR sky130_fd_sc_hd__decap_4
X_5441_ _4598_/X _5441_/Q _4432_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4499__A _4501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_519 VGND VPWR sky130_fd_sc_hd__decap_12
X_5372_ _4743_/X data_out1[2] _4514_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_172_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_530 VGND VPWR sky130_fd_sc_hd__decap_12
X_4323_ _4324_/A _4323_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5099__B1 _5090_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4254_ _4578_/A _4252_/Y _4809_/B _4253_/Y _4254_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_113_287 VGND VPWR sky130_fd_sc_hd__decap_12
X_3205_ _3139_/A _3169_/B _3209_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4185_ _4126_/X _4090_/X _3300_/A _4185_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_68_864 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5123__A _5135_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5422__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_514 VGND VPWR sky130_fd_sc_hd__decap_12
X_3136_ _3073_/C _3096_/B _3136_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_103_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_845 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_867 VGND VPWR sky130_fd_sc_hd__decap_3
X_3067_ _2988_/X _3066_/B _3067_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4962__A _4961_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_761 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5572__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3578__A _3578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_928 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_742 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_405 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4082__A2_N _4081_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_477 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_628 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_263 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_630 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_116 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3969_ _3113_/A _3942_/Y _3969_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5326__B2 _4756_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_357 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_16 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4202__A _4195_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_827 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5017__B _5017_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4856__B _4854_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_950 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_801 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4575__C _4650_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5033__A _5030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_503 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_683 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2863__A2 _2859_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_333 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_193 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4872__A _5547_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4065__A1 _4013_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_761 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_934 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3488__A _3488_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_230 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_764 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_30 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3025__C1 _3024_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_961 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3000__B key_in[47] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_836 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_610 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_493 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_644 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3935__B _3935_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_335 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_655 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_625 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_8 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3654__C _5327_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_904 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_861 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3951__A _3569_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_60 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_714 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_574 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5445__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_639 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_725 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4828__B1 _4819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_224 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3670__B _3669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5556__RESET_B _4295_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4782__A _4700_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_517 VGND VPWR sky130_fd_sc_hd__fill_2
X_4941_ _4642_/A _4847_/X _4531_/X _4940_/X _4941_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3803__B2 _3802_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4872_ _5547_/Q _4838_/B _5548_/Q _4545_/A _4872_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_60_550 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2733__C _2733_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_948 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_3823_ _2914_/X _3822_/X _2914_/X _3822_/X _3823_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4006__B _4007_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3567__B1 _3566_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_3754_ _3725_/Y _3734_/X _3754_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3031__A2 _3030_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_836 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5308__A1 _5264_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_121 VGND VPWR sky130_fd_sc_hd__fill_1
X_2705_ _5299_/A key_in[39] _2705_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_146_655 VGND VPWR sky130_fd_sc_hd__decap_12
X_3685_ _3589_/Y _3683_/X _3727_/A _3685_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__5118__A _5037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4022__A _4014_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5424_ _5424_/D data_out2[22] _4453_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_146_699 VGND VPWR sky130_fd_sc_hd__decap_3
X_5355_ _5355_/A _2698_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_142_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_915 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_819 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_4306_ _4305_/A _4306_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_142_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_937 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_371 VGND VPWR sky130_fd_sc_hd__fill_1
X_5286_ _5256_/A _5285_/X _5286_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_87_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_458 VGND VPWR sky130_fd_sc_hd__fill_1
X_4237_ data_in1[30] _4125_/X _4221_/X _4236_/X _5509_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3384__A1_N _3367_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4168_ _4157_/Y _4168_/B _4168_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_67_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2845__A2 _2842_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_536 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4692__A _5520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3119_ _3077_/A key_in[18] _3119_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5244__B1 _5227_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4099_ _3980_/Y _4098_/X _4099_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_71_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_314 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4598__A2 _4595_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2924__B _2920_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_703 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_714 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5300__B key_in[36] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_764 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_369 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_926 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_414 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_959 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_436 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_419 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_22 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3558__B1 _4661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_600 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2940__A _5497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_611 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_953 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3755__B _3754_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_806 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5333__A2_N _5332_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5028__A _5027_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_614 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_316 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5468__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_349 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_657 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4867__A _4865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_574 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5348__A2_N _5347_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4586__B _4586_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3490__B _3541_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_30 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3089__A2 _3087_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_74 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2836__A2 _2835_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_569 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4038__A1 _4778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2834__B _2795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3246__C1 _3245_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4107__A _4106_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_235 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3946__A _3945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3549__B1 _3533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2850__A _2850_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_970 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_110 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4210__B2 _4209_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_953 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3665__B _3728_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4761__A2 _4757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_452 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_699 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2772__B2 _2771_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3470_ _3499_/A key_in[60] _3470_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5171__C1 _5170_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_701 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3681__A _3681_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5140_ _5133_/Y _5140_/B _5148_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_123_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_533 VGND VPWR sky130_fd_sc_hd__fill_2
X_5071_ _5084_/A _5085_/B _5071_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_96_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_778 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_812 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4816__A3 _4814_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4022_ _4014_/X _4021_/X _4027_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_96_288 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_160 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_620 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5390__RESET_B _4493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_325 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2744__B _5364_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5120__B _5119_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4662__D _4649_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4924_ _5554_/Q _4923_/X _5554_/Q _4923_/X _4924_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4017__A _4775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3252__A2 _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_881 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_892 VGND VPWR sky130_fd_sc_hd__fill_2
X_4855_ _4853_/X _4854_/X _4855_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2760__A _2759_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3806_ _3804_/X _3805_/Y _3806_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_778 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_4786_ _3155_/A _4786_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3004__A2 _3000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_633 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_430 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_964 VGND VPWR sky130_fd_sc_hd__decap_8
X_3737_ _2771_/X _3736_/Y _2771_/X _3736_/Y _3737_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4752__A2 _4745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5493__D _5493_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_934 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_316 VGND VPWR sky130_fd_sc_hd__decap_8
X_3668_ _5346_/X _3667_/X _3668_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_106_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_187 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_967 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_5407_ _5407_/D data_out2[5] _4473_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4687__A _4674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_850 VGND VPWR sky130_fd_sc_hd__decap_4
X_3599_ _3615_/A _3570_/B _5481_/Q _3599_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_88_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3712__B1 _3741_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5338_ _2707_/A key_in[69] _5338_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4837__D _4542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_853 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5478__RESET_B _4388_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_555 VGND VPWR sky130_fd_sc_hd__decap_12
X_5269_ _4636_/A _5265_/X _5266_/X _5267_/X _5268_/X _5270_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_130_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_812 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_981 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5407__RESET_B _4473_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4807__A3 _4802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_322 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2818__A2 _3895_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_491 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_642 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_366 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_472 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_667 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3766__A _3737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_266 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5272__A2_N _5271_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3485__B _3459_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_121 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_20 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4743__A2 _4736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_772 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_176 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_989 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4597__A _4600_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_465 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3703__B1 _5514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_842 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5205__B key_in[65] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_929 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_789 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5210__A2_N _5209_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3006__A _3052_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_333 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_50 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5221__A _4529_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5208__B1 _5303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_910 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_483 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2690__B1 _5365_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5578__D _4263_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_155 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_678 VGND VPWR sky130_fd_sc_hd__decap_6
X_2970_ _2934_/A key_in[78] _2970_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_15_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_82 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3676__A _3676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_728 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_553 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_920 VGND VPWR sky130_fd_sc_hd__fill_2
X_4640_ _4639_/X _4640_/X VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_564 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_931 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_953 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_430 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4195__B1 _4231_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4571_ _5571_/Q _4574_/B _4571_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_129_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_772 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_986 VGND VPWR sky130_fd_sc_hd__fill_2
X_3522_ _4661_/X _3510_/B _3510_/A _3522_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_171_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_809 VGND VPWR sky130_fd_sc_hd__decap_12
X_3453_ _3442_/X _3452_/X _3442_/X _3452_/X _3464_/B VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_143_466 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_628 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4300__A _4303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2739__B _2739_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3384_ _3367_/X _3419_/B _3367_/X _3419_/B _3385_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_842 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5571__RESET_B _4278_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5123_ _5135_/B _5125_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_58_918 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5500__RESET_B _4363_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_428 VGND VPWR sky130_fd_sc_hd__decap_4
X_5054_ _5054_/A _5054_/B _5072_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_111_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_951 VGND VPWR sky130_fd_sc_hd__fill_2
X_4005_ _3958_/X _3984_/X _4007_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_84_269 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2755__A _5301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_815 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3473__A2 key_in[124] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_196 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5488__D _5488_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3690__A2_N _3689_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_37 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4970__A _4958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_177 VGND VPWR sky130_fd_sc_hd__fill_1
X_4907_ _4907_/A _4911_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_21_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_391 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4973__A2 _4971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3586__A _3586_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4838_ _4819_/A _4838_/B _4838_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_166_536 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_227 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_569 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_901 VGND VPWR sky130_fd_sc_hd__fill_2
X_4769_ _4672_/X _4769_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_708 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2736__A1 _2702_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3933__B1 _2989_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_474 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_945 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_45 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_628 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_680 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_520 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_435 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5025__B _5024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5506__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3161__B2 _3160_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_54 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5006__B1_N _5005_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_897 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1002 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_940 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_962 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_269 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_984 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5041__A _5036_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5398__D _4793_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4880__A _4877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_829 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_177 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_497 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_342 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_81 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_525 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3927__C _3926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_558 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4177__B1 _4171_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4716__A2 _4712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_901 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4104__B _4079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_400 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_591 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3943__B _3942_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_617 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4120__A _4114_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_639 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3152__A1 _5013_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_575 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_501 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_597 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_225 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_166 VGND VPWR sky130_fd_sc_hd__decap_8
X_2953_ _2930_/Y _2988_/B _2953_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2884_ _2733_/A _2884_/B _5523_/Q _2884_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_31_895 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2805__A2_N _2804_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4623_ _2861_/A _3077_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_260 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3915__B1 _3058_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4554_ _4554_/A _4547_/B _4554_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4949__B _4949_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3853__B _3852_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3505_ _5143_/X _3504_/X _5143_/A _3504_/X _3505_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5529__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4485_ _4483_/X _4485_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_403 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5126__A _5125_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_274 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4030__A _3905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_3436_ _3436_/A _3436_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_650 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_715 VGND VPWR sky130_fd_sc_hd__decap_4
X_3367_ _3321_/Y _3349_/A _4661_/X _3367_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4965__A _4554_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1005 VGND VPWR sky130_fd_sc_hd__decap_12
X_5106_ _5134_/A _5124_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_383 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_171 VGND VPWR sky130_fd_sc_hd__fill_2
X_3298_ _3268_/Y _3271_/X _3267_/Y _3298_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_57_258 VGND VPWR sky130_fd_sc_hd__decap_12
X_5037_ _4975_/X _5037_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_73_718 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_450 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3446__A2 key_in[123] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_910 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_770 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_612 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4643__B2 _4616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2932__B key_in[45] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4205__A _4126_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2709__A1 _4636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3906__B1 _5523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2709__B2 _2708_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_720 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5493__RESET_B _4371_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3763__B _3761_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3382__B2 _3381_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_455 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5036__A _5468_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5422__RESET_B _4456_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_733 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3134__A1 _3133_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4875__A _4876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_777 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_661 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3685__A2 _3683_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_726 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_694 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4594__B _4590_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_247 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_472 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_217 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_526 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4634__B2 _4616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1012 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_604 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_51 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3938__B _3937_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2842__B _2842_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_800 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_84 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2948__A1 _4661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_161 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4115__A _4115_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_169 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_670 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_183 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_844 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_194 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3535__A2_N _3534_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3954__A _3904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_399 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_731 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5362__A2 _5361_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3673__B _3651_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3373__B2 _3372_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_701 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_403 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_4270_ _4271_/A _4270_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_147 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3125__A1 _4996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_255 VGND VPWR sky130_fd_sc_hd__decap_12
X_3221_ _3145_/X _3291_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3092__A1_N _3937_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_288 VGND VPWR sky130_fd_sc_hd__decap_6
X_3152_ _5013_/A _3195_/B _3196_/B _3197_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_67_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_206 VGND VPWR sky130_fd_sc_hd__decap_8
X_3083_ _3128_/A _3057_/Y _3048_/Y _3083_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3428__A2 _3427_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4009__B _4008_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_987 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_946 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_445 VGND VPWR sky130_fd_sc_hd__decap_12
X_3985_ _3958_/X _3962_/X _3957_/X _3985_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_22_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4670__D _4669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2939__B2 _2938_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2936_ _4637_/X _2932_/X _2933_/X _2934_/X _2935_/X _2936_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_50_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_2867_ _3902_/C _3032_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3864__A _3843_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1001 VGND VPWR sky130_fd_sc_hd__decap_12
X_4606_ _4605_/X _4609_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_731 VGND VPWR sky130_fd_sc_hd__fill_1
X_2798_ _3671_/A _3870_/A _5327_/A _2961_/A _2799_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3583__B _3570_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_753 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_4537_ _4893_/A _4537_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_172_881 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_4468_ _4468_/A _4468_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_136 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_233 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_158 VGND VPWR sky130_fd_sc_hd__fill_1
X_3419_ _3419_/A _3419_/B _3419_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_113_970 VGND VPWR sky130_fd_sc_hd__fill_2
X_4399_ _4402_/A _4399_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_821 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2927__B _2925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2875__B1 _2857_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3104__A _2885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_932 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_420 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_913 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2943__A _2943_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_clock clkbuf_4_9_0_clock/A _5372_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_626 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__A2 _4847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_21 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_32 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_333 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_681 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_815 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_303 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_185 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_836 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_859 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_858 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4589__B _4588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__B _3364_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3355__A1 _3287_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_550 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3924__D _3923_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_520 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_745 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_810 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_439 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2866__B1 _2858_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_589 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3014__A _3014_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_846 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_740 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_442 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3949__A _4664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_976 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_902 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_773 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3668__B _3667_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_732 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_445 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5374__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_776 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_618 VGND VPWR sky130_fd_sc_hd__decap_12
X_3770_ _4707_/A _3770_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_13_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_692 VGND VPWR sky130_fd_sc_hd__decap_4
X_2721_ _2713_/X _2720_/X _2713_/X _2720_/X _2722_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_815 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3594__B2 _3593_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_837 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3684__A _3589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5440_ _4593_/Y _5440_/Q _4434_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_66_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_807 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_5371_ _5371_/D data_out1[1] _4515_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_126_572 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_199 VGND VPWR sky130_fd_sc_hd__decap_12
X_4322_ _4324_/A _4322_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_891 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_542 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5099__A1 _4896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5099__B2 _4806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_607 VGND VPWR sky130_fd_sc_hd__decap_3
X_4253_ _4524_/A _4629_/D _4519_/X _4253_/D _4253_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_99_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_299 VGND VPWR sky130_fd_sc_hd__decap_6
X_3204_ _3175_/Y _3203_/B _3217_/A _3213_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_68_843 VGND VPWR sky130_fd_sc_hd__decap_8
X_4184_ data_in1[27] _4125_/X _4167_/X _4183_/Y _5506_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_79_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_707 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_718 VGND VPWR sky130_fd_sc_hd__decap_12
X_3135_ _3069_/A _3099_/B _3068_/Y _3135_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_67_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_898 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_824 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_984 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_526 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_228 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_3066_ _2991_/B _3066_/B _3066_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_82_345 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4962__B _4960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5271__A1 _4827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2763__A _2686_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_570 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3282__B1 _3353_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_890 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3578__B _3575_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_417 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5496__D _5496_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_242 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_428 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3034__B1 _3033_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3968_ _3925_/A _3945_/B _3924_/Y _3968_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_137_804 VGND VPWR sky130_fd_sc_hd__fill_2
X_2919_ _2918_/A _2918_/B _2930_/A _2925_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_136_303 VGND VPWR sky130_fd_sc_hd__decap_12
X_3899_ _3883_/Y _3921_/B _3899_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_137_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_185 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_678 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_306 VGND VPWR sky130_fd_sc_hd__decap_8
X_5569_ _5569_/D _5569_/Q _4280_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4202__B _4232_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_715 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5314__A _5284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_832 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2848__B1 _2806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5033__B _5032_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_695 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2863__A3 _2860_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_857 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4872__B _4838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_345 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5397__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4065__A2 _4064_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3769__A _2842_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_732 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_592 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3488__B _3488_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_406 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_776 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_53 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3025__B1 _2996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_86 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_804 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4773__B1 data_out1[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_314 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_655 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_677 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_572 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3505__A1_N _5143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_704 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_938 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_72 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4828__A1 _4541_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5224__A _5252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_353 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_813 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_846 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_131 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_805 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3679__A _3615_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_153 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_687 VGND VPWR sky130_fd_sc_hd__decap_12
X_4940_ _4918_/A _4938_/Y _4949_/B _4940_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3264__B1 _3222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_220 VGND VPWR sky130_fd_sc_hd__fill_2
X_4871_ _4871_/A _4876_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_21_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_776 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5525__RESET_B _4332_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3822_ _3818_/X _3821_/Y _3822_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_159_940 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3016__B1 _3036_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_951 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_595 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3567__A1 _3564_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3753_ _3636_/Y _3751_/X _3752_/X _3753_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_20_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4764__B1 data_out1[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_483 VGND VPWR sky130_fd_sc_hd__decap_12
X_2704_ _2687_/X _2688_/X _2686_/Y _2704_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_118_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_848 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4303__A _4303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5308__A2 _5307_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3684_ _3589_/Y _3683_/X _3727_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_145_133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_667 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_604 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5118__B _5129_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5423_ _4719_/X data_out2[21] _4454_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_118_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_615 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4022__B _4021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_5354_ data_in2[5] _5222_/X _5321_/X _5353_/X _5354_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_99_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_242 VGND VPWR sky130_fd_sc_hd__fill_2
X_4305_ _4305_/A _4305_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_873 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3351__A2_N _3365_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_350 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_5285_ _5256_/B _5275_/B _5285_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_895 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5134__A _5134_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_225 VGND VPWR sky130_fd_sc_hd__decap_3
X_4236_ _3676_/A _4236_/B _4236_/C _4236_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5026__A1_N _5563_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_4167_ _4126_/X _4090_/X _4791_/X _4167_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_55_312 VGND VPWR sky130_fd_sc_hd__fill_2
X_3118_ _3043_/X key_in[50] _3118_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_643 VGND VPWR sky130_fd_sc_hd__fill_2
X_4098_ _3175_/Y _5540_/Q _3175_/A _4097_/Y _4098_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3589__A _5517_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5244__B2 _5243_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_827 VGND VPWR sky130_fd_sc_hd__decap_4
X_3049_ _5463_/Q _3047_/B _3048_/Y _3128_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3255__B1 _3254_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2924__C _2924_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_890 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_743 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_938 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3007__B1 _3006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4204__C1 _4203_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_45 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3558__A1 _3522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4755__B1 data_out1[9] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_921 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_971 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5309__A _5306_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_494 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4213__A _4794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_475 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_626 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_636 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4867__B _4866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_586 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5044__A _5056_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_556 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_971 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3494__B1 _3465_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_183 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_559 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4038__A2 _4036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3499__A _3499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_838 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_315 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3246__B1 _3216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4994__B1 _4993_/Y VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_clock clkbuf_3_6_0_clock/A clkbuf_3_6_0_clock/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_14_264 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_40 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_91 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3549__A1 _5154_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3549__B2 _3534_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3946__B _3945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2850__B _2850_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_910 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_84 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5219__A _5281_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4123__A _4092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5412__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_964 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_317 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3962__A _3959_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_328 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_840 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5171__B1 _4542_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3681__B _3680_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_404 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_884 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5562__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_501 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4081__A2_N _4080_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_692 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_394 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_691 VGND VPWR sky130_fd_sc_hd__decap_8
X_5070_ _5068_/A _5067_/X _5085_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_85_908 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_556 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_267 VGND VPWR sky130_fd_sc_hd__decap_8
X_4021_ _4016_/X _4020_/Y _4021_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_65_632 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_805 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_816 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_602 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3237__B1 _3257_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_849 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_337 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2744__C _2744_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4923_ _4921_/X _4922_/X _4923_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4017__B _3990_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4854_ _4840_/X _4844_/X _4854_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_33_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_370 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_707 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_770 VGND VPWR sky130_fd_sc_hd__fill_2
X_3805_ _3804_/A _3803_/X _3805_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_119_601 VGND VPWR sky130_fd_sc_hd__fill_2
X_4785_ _4784_/X _4781_/X data_out1[23] _4782_/X _4785_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_20_256 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3004__A3 _3001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5129__A _5129_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3736_ _3726_/Y _3733_/X _3735_/Y _3736_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_118_122 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_645 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4034__A2_N _4033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_442 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_290 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_829 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_166 VGND VPWR sky130_fd_sc_hd__decap_6
X_3667_ _3666_/X _3667_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4968__A _3052_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_114 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3872__A _3871_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5406_ _5406_/D data_out2[4] _4474_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_133_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5162__B1 _5160_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_979 VGND VPWR sky130_fd_sc_hd__decap_4
X_3598_ data_in1[1] _3581_/X _3583_/X _3597_/X _3598_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3712__A1 _2717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_713 VGND VPWR sky130_fd_sc_hd__fill_2
X_5337_ _2707_/A key_in[5] _5337_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_681 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_383 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_245 VGND VPWR sky130_fd_sc_hd__decap_3
X_5268_ _5234_/A key_in[99] _5303_/A _5268_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_130_865 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_960 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_4219_ _4092_/X _4219_/B _4218_/X _4219_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_5199_ _5480_/Q _5199_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_18_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_45 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_451 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5447__RESET_B _4425_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_326 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3112__A _3038_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_501 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4976__B1 _4975_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_534 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5435__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_735 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_910 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_227 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5039__A _5037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_954 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_976 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_924 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4878__A _4863_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_475 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_400 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_637 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3782__A _3743_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5153__B1 _5146_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_840 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_478 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3703__A1 _5253_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_629 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3703__B2 _2918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_74 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3006__B _3052_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3467__B1 _3466_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5208__A1 _5234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4112__A1_N _4786_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_922 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4118__A _4016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_495 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3022__A _2997_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2690__B2 _2689_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_646 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4967__B1 _4555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_90 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_562 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3957__A _3133_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2861__A _2861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_532 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3676__B _3674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4719__B1 data_out2[21] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4195__A1 _3466_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4570_ _5129_/A _4574_/B _5570_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_156_751 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3383__A1_N _3373_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_750 VGND VPWR sky130_fd_sc_hd__decap_12
X_3521_ _3520_/Y _3521_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4788__A _3178_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3692__A _3671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_282 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_231 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5144__B1 _5052_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3452_ _3452_/A _3452_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_489 VGND VPWR sky130_fd_sc_hd__fill_2
X_3383_ _3373_/X _3382_/X _3373_/X _3382_/X _3419_/B VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_97_510 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_821 VGND VPWR sky130_fd_sc_hd__decap_3
X_5122_ _5122_/A _5138_/A _5135_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_5053_ _5065_/A _5052_/X _5065_/A _5052_/X _5054_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_289 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_930 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_749 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_941 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_397 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_248 VGND VPWR sky130_fd_sc_hd__decap_3
X_4004_ _3957_/X _3982_/X _4008_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_37_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2755__B key_in[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_473 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5540__RESET_B _4314_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_635 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5458__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_977 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4970__B _4962_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_871 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3867__A _3823_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4906_ _4896_/X _4903_/Y _4904_/X _4905_/Y _4806_/X _4906_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XANTENNA__5347__A2_N _5346_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4973__A3 _4972_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3039__B1_N _3038_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4837_ _5543_/Q _4837_/B _4541_/A _4542_/A _4838_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_21_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_576 VGND VPWR sky130_fd_sc_hd__fill_2
X_4768_ _3895_/A _4757_/X data_out1[15] _4758_/X _4768_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_135_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_924 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3933__A1 _3721_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2736__A2 _2722_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3933__B2 _3932_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4698__A _4672_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3719_ _3765_/A _3679_/B _5261_/A _3719_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_119_486 VGND VPWR sky130_fd_sc_hd__fill_2
X_4699_ _4699_/A _4699_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_434 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_754 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_905 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_927 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3107__A _3060_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_692 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_447 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_386 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5322__A _5322_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_805 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_142 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5041__B _5040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_76 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4880__B _4878_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_860 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_871 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_487 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_893 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_343 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_504 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_503 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_42 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4177__B2 _4176_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_751 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4104__C _4055_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_913 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_412 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4401__A _4402_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_927 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4120__B _4120_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_128 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_285 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_692 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_296 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3152__A2 _3195_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_554 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_684 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2856__A _2814_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_952 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_741 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_465 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3687__A _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2952_ _2930_/Y _2988_/B _2952_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_96_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_392 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A clkbuf_3_6_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_2883_ _5355_/A _2884_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_4622_ _2934_/A _2861_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_30_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_570 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3915__B2 _3914_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4553_ _4553_/A _4547_/B _4553_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_156_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_743 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_220 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_754 VGND VPWR sky130_fd_sc_hd__decap_8
X_3504_ _4640_/X _3500_/X _3501_/X _3502_/X _3503_/X _3504_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4311__A _4304_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4484_ _4483_/X _4484_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_467 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_562 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5126__B _5124_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_415 VGND VPWR sky130_fd_sc_hd__decap_12
X_3435_ _3435_/A _3432_/B _3459_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4030__B _4028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4634__A1_N _4616_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3366_ _3366_/A _3362_/B _3388_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4965__B _4955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_662 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_727 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_513 VGND VPWR sky130_fd_sc_hd__fill_2
X_5105_ _5104_/X _5134_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2766__A _2766_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1017 VGND VPWR sky130_fd_sc_hd__decap_3
X_3297_ _5470_/Q _3295_/X _3296_/X _3297_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_57_226 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_941 VGND VPWR sky130_fd_sc_hd__fill_2
X_5036_ _5468_/Q _5036_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_39_963 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5499__D _5499_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_782 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_484 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_933 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4981__A _4982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_590 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_808 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_156 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_465 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3597__A _3579_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_329 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_638 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_515 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_846 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_351 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4205__B _4090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_323 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_559 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3906__A1 _2918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2709__A2 _2705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_401 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_924 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3906__B2 _3905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_539 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5317__A _5317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4221__A _4126_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3763__C _3762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_467 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_713 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_724 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_clock clkbuf_4_5_0_clock/A _5413_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_135_798 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_949 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_768 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3134__A2 _3133_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4875__B _4874_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_960 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_502 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_77 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_738 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5462__RESET_B _4408_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_492 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5052__A _5052_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5239__A2_N _5238_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_42 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4891__A _4891_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_495 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_432 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_999 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_262 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_189 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3300__A _3300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_137 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_813 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2948__A2 _2916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_151 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_812 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_162 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4115__B _4115_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_823 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_173 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_323 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_682 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_195 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5347__B1 _5333_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_304 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_366 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3954__B _3953_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_581 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5227__A _5256_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_253 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4858__C1 _4857_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_768 VGND VPWR sky130_fd_sc_hd__fill_2
X_3220_ _3148_/A key_in[85] _3220_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3125__A2 _3122_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_779 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_960 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_204 VGND VPWR sky130_fd_sc_hd__fill_1
X_3151_ _5013_/A _3195_/B _3196_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_94_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3082_ _4985_/X _3081_/B _3127_/B _3128_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_82_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_936 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4306__A _4305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3210__A _3207_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3984_ _3982_/X _3983_/Y _3984_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_813 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_2935_ _2968_/A key_in[109] _2828_/X _2935_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_148_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3061__A1 _3060_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_879 VGND VPWR sky130_fd_sc_hd__decap_12
X_2866_ _2858_/Y _2865_/X _2858_/Y _2865_/X _3801_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_838 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3864__B _3862_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4605_ _4646_/A _4605_/B _4605_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_11_1013 VGND VPWR sky130_fd_sc_hd__decap_6
X_2797_ _2797_/A _2961_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5137__A _5108_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4041__A _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3583__C _3583_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4536_ _4529_/X _4893_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_105_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_562 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_893 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_735 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_48 VGND VPWR sky130_fd_sc_hd__decap_4
X_4467_ _4468_/A _4467_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3880__A _3835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_256 VGND VPWR sky130_fd_sc_hd__fill_2
X_3418_ _3403_/X _3417_/X _3403_/X _3417_/X _3436_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4398_ _4402_/A _4398_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_289 VGND VPWR sky130_fd_sc_hd__fill_2
X_3349_ _3349_/A _3419_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_470 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_535 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2875__B2 _2887_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2927__C _2926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_354 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_900 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_505 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_527 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_782 VGND VPWR sky130_fd_sc_hd__fill_2
X_5019_ _5002_/Y _5019_/B _5019_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_27_955 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_432 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_605 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2943__B _2943_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_796 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_947 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4216__A _4231_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3120__A _3077_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4214__B1_N _4213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_800 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_643 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_827 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_315 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2866__A2_N _2865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4001__B1 _5527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5047__A _5047_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_808 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3493__C _3493_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3355__A2 _3309_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_893 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3790__A _3765_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_768 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_535 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2866__B2 _2865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_825 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3014__B _3014_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_858 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_454 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5519__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_711 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_498 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4126__A _4537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_593 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3030__A _3030_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_621 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4240__B1 _3848_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2720_ _2744_/C _2719_/X _2744_/C _2719_/X _2720_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_676 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3684__B _3683_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_156 VGND VPWR sky130_fd_sc_hd__decap_12
X_5370_ _4740_/X data_out1[0] _4516_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5384__RESET_B _4500_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4321_ _4324_/A _4321_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5099__A2 _5097_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_234 VGND VPWR sky130_fd_sc_hd__fill_2
X_4252_ _4576_/X _4252_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_822 VGND VPWR sky130_fd_sc_hd__fill_2
X_3203_ _3175_/Y _3203_/B _3217_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_4183_ _4092_/X _4183_/B _4183_/C _4183_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_67_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_941 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3205__A _3139_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3134_ _3133_/A _3133_/B _3144_/A _3139_/A VGND VPWR sky130_fd_sc_hd__a21o_4
Xclkbuf_0_clock clock clkbuf_0_clock/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_83_836 VGND VPWR sky130_fd_sc_hd__fill_2
X_3065_ _3065_/A _3065_/B _3066_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_103_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_195 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5271__A2 _5270_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2763__B _2711_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3282__A1 _3211_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_947 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_733 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_766 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_608 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3034__A1 _3032_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3967_ _3110_/A _3965_/X _3966_/Y _3972_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_50_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3875__A _3875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_991 VGND VPWR sky130_fd_sc_hd__decap_12
X_2918_ _2918_/A _2918_/B _2930_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xclkbuf_1_0_0_clock clkbuf_0_clock/X clkbuf_2_1_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_109_507 VGND VPWR sky130_fd_sc_hd__fill_2
X_3898_ _3883_/Y _3921_/B _3898_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_109_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_613 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2793__B1 _2790_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_47 VGND VPWR sky130_fd_sc_hd__decap_4
X_2849_ _2849_/A _2849_/B _2850_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_148_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_5568_ _4567_/X _5568_/Q _4281_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_151_318 VGND VPWR sky130_fd_sc_hd__decap_6
X_4519_ _4518_/X _4519_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5499_ _5499_/D _3010_/A _4364_/X _5430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_120_727 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5314__B _5313_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_598 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2848__A1 _2784_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3115__A _3112_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_814 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2954__A _2927_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_495 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4872__C _5548_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_56 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_357 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5330__A _5330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_903 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_880 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_435 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_744 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3488__C _3488_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_43 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3025__A1 data_in2[15] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4222__B1 _4212_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3785__A _3831_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_287 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3091__A1_N _3112_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4773__A1 _3113_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4773__B2 _4770_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_326 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_674 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_634 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_871 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_318 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_689 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_608 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_clock clkbuf_3_2_0_clock/A clkbuf_4_5_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_97_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_416 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4828__A2 _4818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5224__B _5252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_215 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2839__A1 _2838_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_790 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_641 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5040__A2_N _5039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_302 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_61 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2864__A _2907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3679__B _3679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_817 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3264__A1 _3291_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3992__B1_N _4018_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_722 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_4870_ _4857_/A _4870_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_243 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5491__CLK _5430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3821_ _3799_/B _3819_/Y _3820_/Y _3821_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_21_928 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_276 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3016__B2 _3015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3059__A1_N _3039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3695__A _3676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_963 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4764__A1 _3875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3567__A2 _3565_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3752_ _3636_/Y _3751_/X _3752_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3689__A1_N _2689_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4764__B2 _4758_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_996 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2775__B1 _2784_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2703_ _5358_/A _2702_/X _2722_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__5565__RESET_B _4285_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_495 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_483 VGND VPWR sky130_fd_sc_hd__decap_4
X_3683_ _3603_/A _2876_/A _5513_/Q _3682_/Y _3683_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_145 VGND VPWR sky130_fd_sc_hd__decap_12
X_5422_ _5422_/D data_out2[20] _4456_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_127_893 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_690 VGND VPWR sky130_fd_sc_hd__decap_8
X_5353_ _2696_/A _5351_/X _5352_/Y _5353_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_99_232 VGND VPWR sky130_fd_sc_hd__decap_4
X_4304_ _4304_/A _4305_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_405 VGND VPWR sky130_fd_sc_hd__decap_12
X_5284_ _5515_/Q _5284_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_114_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_727 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5134__B _5122_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_395 VGND VPWR sky130_fd_sc_hd__fill_2
X_4235_ _4229_/X _4234_/B _4236_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_68_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_803 VGND VPWR sky130_fd_sc_hd__decap_8
X_4166_ data_in1[26] _4125_/X _4144_/X _4165_/Y _4166_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_56_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_685 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_471 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_482 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2774__A _2735_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3117_ _3116_/A _3115_/X _3116_/X _3131_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_67_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_4097_ _5540_/Q _4097_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5150__A _5147_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_357 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_3048_ _3048_/A _3048_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_130_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3255__A1 _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_305 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_688 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2924__D _2923_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_210 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_593 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_221 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_530 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_755 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_215 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3007__A1 _5462_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4204__B1 _4185_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4999_ _4559_/A _4998_/X _4559_/A _4998_/X _4999_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4755__A1 _3759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3558__A2 _3536_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_911 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4755__B2 _4746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5309__B _5308_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_432 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4213__B _4212_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_966 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_648 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_125 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5325__A _5325_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_874 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_928 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5044__B _5057_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3494__A1 _3465_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_994 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4691__B1 data_out2[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5060__A _5072_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3246__A1 data_in2[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_327 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_64 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_75 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_349 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4994__A1 _4896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_97 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4994__B2 _4806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_30 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4404__A _4267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3549__A2 _3532_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_52 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_760 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3411__A2_N _3410_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2757__B1 _2828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_270 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5219__B _5217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4123__B _4123_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_471 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_668 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_808 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_988 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_167 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_475 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3962__B _3961_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_126 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5171__A1 _5478_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2859__A _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_852 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5235__A _5236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_681 VGND VPWR sky130_fd_sc_hd__decap_8
X_4020_ _4020_/A _4018_/X _4019_/Y _4020_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_111_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_983 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_460 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4682__B1 data_out2[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_920 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_644 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3237__B2 _3236_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4910__A1_N _5553_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4922_ _5553_/Q _4908_/X _4922_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4853_ _4852_/A _4851_/X _4852_/X _4853_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_60_382 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_719 VGND VPWR sky130_fd_sc_hd__decap_12
X_3804_ _3804_/A _3803_/X _3804_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4314__A _4312_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4784_ _3108_/A _4784_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_268 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5129__B _5129_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3735_ _3734_/X _3735_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_119_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_988 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_402 VGND VPWR sky130_fd_sc_hd__fill_2
X_3666_ _3666_/A _3666_/B _3666_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4968__B _4968_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_947 VGND VPWR sky130_fd_sc_hd__decap_4
X_5405_ _4682_/X data_out2[3] _4475_/X _5402_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5387__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5162__A1 _5154_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2769__A _2769_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3597_ _3579_/A _3595_/X _3596_/Y _3597_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_88_703 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3712__A2 _3710_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5336_ _5299_/A key_in[37] _5336_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_5267_ _5236_/A key_in[67] _5267_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_19 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_877 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_972 VGND VPWR sky130_fd_sc_hd__decap_4
X_4218_ _4215_/Y _4218_/B _4218_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_102_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3476__A1 _5116_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5198_ _5198_/A _5198_/B _5198_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_4149_ _4147_/X _4149_/B _4173_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_141_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_36 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_508 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_496 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_891 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_338 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3112__B _3112_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_135 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4976__A1 _4555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_23 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2987__B1 _3064_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_168 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5487__RESET_B _4378_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_546 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_708 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5416__RESET_B _4463_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_729 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_270 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5039__B _5038_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_730 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3400__A1 _3396_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_988 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_66 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_785 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_936 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4878__B _4868_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_412 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_935 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3782__B _3782_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_649 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5153__A1 _5133_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5153__B2 _5152_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_852 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3164__B1 _3107_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_456 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_863 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3703__A2 _5523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_373 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4894__A _4656_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_769 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3467__A1 _4786_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_931 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_942 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_964 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_290 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3303__A _3108_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_817 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5208__A2 key_in[97] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2713__A1_N _2704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_379 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4118__B _4119_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_945 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3022__B _3065_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4967__B2 _4966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_872 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3957__B _3956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2978__B1 _2977_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_883 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2861__B key_in[75] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3676__C _3675_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4134__A _4101_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4719__A1 _4718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4719__B2 _4713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4109__A2_N _4108_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4195__A2 _4193_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3973__A _3972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_977 VGND VPWR sky130_fd_sc_hd__decap_6
X_3520_ _5541_/Q _3520_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_116_605 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_999 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_762 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_947 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3692__B _3674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_958 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5144__A1 _5571_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_272 VGND VPWR sky130_fd_sc_hd__decap_3
X_3451_ _3450_/A _3449_/Y _3450_/X _3452_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_109_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_243 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_3382_ _3414_/B _3381_/Y _3414_/B _3381_/Y _3382_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_991 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_522 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2902__B1 _2900_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5121_ _5121_/A _5119_/X _5138_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_69_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_866 VGND VPWR sky130_fd_sc_hd__decap_4
X_5052_ _5052_/A _5051_/X _5052_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_57_419 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_611 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_780 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_110 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_633 VGND VPWR sky130_fd_sc_hd__decap_3
X_4003_ _3175_/Y _4001_/X _4002_/X _4003_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__4309__A _4305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_132 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3213__A _3213_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_603 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_794 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_124 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_647 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_349 VGND VPWR sky130_fd_sc_hd__fill_2
X_4905_ _4900_/A _4905_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3867__B _3847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_691 VGND VPWR sky130_fd_sc_hd__fill_2
X_4836_ _4836_/A _4840_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4044__A _4011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_190 VGND VPWR sky130_fd_sc_hd__fill_2
X_4767_ _5494_/Q _3895_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3883__A _3871_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3933__A2 _4720_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3718_ data_in1[7] _3697_/X _3699_/X _3717_/Y _3718_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_4_209 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_722 VGND VPWR sky130_fd_sc_hd__decap_12
X_4698_ _4672_/X _4699_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_161_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_3649_ _3626_/X _3631_/B _3649_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_136_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_298 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3107__B _3107_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5319_ _5281_/A _5319_/B _5319_/C _5319_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_103_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_23 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_459 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3449__A1 _5473_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_57 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4219__A _4092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_452 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3123__A _4996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5402__CLK _5402_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_997 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_839 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_967 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_809 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_1_0_clock clkbuf_4_1_0_clock/A _5429_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_71_455 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_321 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5552__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_544 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_853 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_577 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_897 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4889__A _4886_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3793__A _3767_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_560 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_571 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_732 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_457 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_231 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3137__B1 _3136_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_308 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_253 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_500 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3688__A1 _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4120__C _4118_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_630 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_566 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_717 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2856__B _2840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_931 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_290 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4129__A _4128_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3033__A _3090_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_452 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4033__A2_N _4032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_474 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_636 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3968__A _3925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_422 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_433 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_444 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2872__A _2872_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_989 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3687__B _3686_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2951_ _2989_/A _2989_/B _2950_/X _2988_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_16_894 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_864 VGND VPWR sky130_fd_sc_hd__decap_12
X_2882_ data_in2[11] _2731_/X _2854_/X _2881_/Y _2882_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_89_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_886 VGND VPWR sky130_fd_sc_hd__fill_2
X_4621_ _5301_/A _2934_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5365__A1 _5364_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4799__A _5543_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_925 VGND VPWR sky130_fd_sc_hd__fill_2
X_4552_ _4944_/A _4547_/B _4552_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_156_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_3503_ _3528_/A key_in[125] _3408_/X _3503_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_143_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_4483_ _4469_/A _4483_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3208__A _3144_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_479 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_265 VGND VPWR sky130_fd_sc_hd__decap_6
X_3434_ _3519_/A _3364_/B _4731_/X _3434_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_98_842 VGND VPWR sky130_fd_sc_hd__decap_12
X_3365_ _3316_/C _3365_/B _3366_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_5104_ _5104_/A _5103_/X _5104_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5425__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_674 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_162 VGND VPWR sky130_fd_sc_hd__fill_2
X_3296_ _5470_/Q _3295_/X _3296_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2938__B1_N _2937_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5035_ _4870_/X _5033_/X _5034_/X _5023_/A _4930_/X _5035_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4039__A _4039_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_986 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_923 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_720 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_580 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4981__B _4980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3878__A _3873_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5575__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_135 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5053__B1 _5065_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3597__B _3595_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_831 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_803 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_842 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_505 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_302 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2811__C1 _2810_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_527 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4205__C _4794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_538 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_869 VGND VPWR sky130_fd_sc_hd__decap_12
X_4819_ _4819_/A _4818_/X _4819_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3367__B1 _4661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3906__A2 _3905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4502__A _4501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2709__A3 _2706_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_413 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_947 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5317__B _5317_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_958 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4221__B _3569_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_552 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3118__A _3043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_928 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_479 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3825__A2_N _3824_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_736 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_853 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2957__A _5223_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_875 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5052__B _5051_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_547 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_452 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3382__A1_N _3414_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_54 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_517 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_463 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4891__B _4889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_282 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3788__A _3788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_444 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5431__RESET_B _4444_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_904 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_959 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_842 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_141 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_302 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_173 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_185 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5347__B2 _5346_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_560 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4412__A _4419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_378 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5227__B _5227_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_541 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_232 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3028__A _2999_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5448__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_265 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_939 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4858__B1 _4531_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_747 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_438 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2867__A _3902_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3965__A1_N _3954_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5346__A2_N _5345_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3150_ _4638_/X _3146_/X _3147_/X _3148_/X _3149_/X _3195_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_94_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_823 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_845 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_333 VGND VPWR sky130_fd_sc_hd__decap_3
X_3081_ _5464_/Q _3081_/B _3127_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5519__RESET_B _4339_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_411 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_934 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_956 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3698__A _4537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_591 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_904 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5035__B1 _5023_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_3983_ _3858_/Y _3981_/X _3983_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3210__B _3210_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2934_ _2934_/A key_in[77] _2934_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3061__A2 _3060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_2865_ _2907_/A _2863_/X _2864_/X _2865_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_148_357 VGND VPWR sky130_fd_sc_hd__fill_2
X_4604_ _5443_/Q _4601_/B _4603_/Y _5443_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_163_316 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3864__C _3863_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4322__A _4324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4010__A1 _4003_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2796_ _2785_/Y _2795_/X _2785_/Y _2795_/X _2796_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_733 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5137__B _5137_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4535_ _5543_/Q _4542_/B _5543_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_850 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4041__B _4041_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_703 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_27 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_939 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_38 VGND VPWR sky130_fd_sc_hd__decap_4
X_4466_ _4468_/A _4466_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_213 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_747 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3880__B _3878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_769 VGND VPWR sky130_fd_sc_hd__fill_2
X_3417_ _3416_/A _3415_/Y _3416_/X _3417_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_113_950 VGND VPWR sky130_fd_sc_hd__fill_2
X_4397_ _4397_/A _4402_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_3348_ _3333_/Y _3347_/X _3333_/Y _3347_/X _3349_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_611 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_845 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_622 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_482 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4992__A _4992_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_3279_ _3213_/A _3244_/B _3356_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_5018_ _5017_/A _5017_/B _5017_/X _5021_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_73_539 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2800__B1_N _2799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_550 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5026__B1 _5563_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_403 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4216__B _4203_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_594 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3120__B key_in[82] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_611 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_650 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_970 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_812 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_655 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_805 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5328__A _5327_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_839 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4232__A _4195_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4001__A1 _3062_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_327 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4001__B2 _4000_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5047__B _5045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_210 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_755 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_563 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_371 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_585 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3790__B _3679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_609 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_823 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_460 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_599 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_994 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_525 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_528 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_336 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_967 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4407__A _4411_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3311__A _3312_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_285 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4240__A1 _4222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_789 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_992 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_491 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_688 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4142__A _4092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_541 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_703 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3751__B1 _5321_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3274__A1_N _3250_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4320_ _4324_/A _4320_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_585 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_436 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5099__A3 _5098_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4251_ _4517_/Y _4668_/Y _4255_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3503__B1 _3408_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3202_ _3177_/Y _3201_/X _3177_/Y _3201_/X _3203_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4182_ _4168_/Y _4182_/B _4183_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_68_834 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1007 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3205__B _3169_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3133_ _3133_/A _3133_/B _3144_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_94_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_804 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_697 VGND VPWR sky130_fd_sc_hd__fill_2
X_3064_ _3064_/A _3020_/Y _3064_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_36_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_369 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4317__A _4312_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3221__A _3145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3282__A2 _3356_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_909 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_778 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3966_ _3110_/A _3965_/X _3966_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3034__A2 _3032_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_121 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3875__B _3850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_655 VGND VPWR sky130_fd_sc_hd__fill_2
X_2917_ _2888_/Y _2916_/Y _2888_/Y _2916_/Y _2918_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3897_ _3895_/X _3896_/Y _3921_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_148_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5148__A _5132_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2793__A1 _4637_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3990__B1 _3987_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2793__B2 _2792_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2848_ _2784_/A _2847_/X _2806_/X _2849_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_136_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_135 VGND VPWR sky130_fd_sc_hd__decap_4
X_5567_ _4566_/X _4566_/A _4282_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4987__A _4987_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_541 VGND VPWR sky130_fd_sc_hd__fill_2
X_2779_ _2778_/X _2779_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3891__A _3890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_307 VGND VPWR sky130_fd_sc_hd__fill_2
X_4518_ _4518_/A _4518_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_382 VGND VPWR sky130_fd_sc_hd__fill_2
X_5498_ _5498_/D _2959_/A _4365_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4449_ _4449_/A _4449_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_886 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_812 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2848__A2 _2847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_845 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3115__B _3115_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_889 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_366 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_377 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_13 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2954__B _2952_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4872__D _4545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_89 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_509 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3131__A _3131_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_403 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3488__D _3487_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_756 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2970__A _2934_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3025__A2 _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4222__A1 _3848_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_953 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3785__B _3785_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4773__A2 _4769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_299 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_474 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3981__B1 _3020_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_625 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_636 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_647 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4897__A _5456_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_617 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_680 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_894 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_178 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_566 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_428 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5224__C _5513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2839__A2 _2837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_290 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5238__B1 _5236_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_826 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_314 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2864__B _2863_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3679__C _4750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3264__A2 key_in[118] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3041__A _2861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_572 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_881 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_285 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_520 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_907 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3976__A _4533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2880__A _2855_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3820_ _3773_/X _3820_/B _3774_/X _3820_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_32_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_575 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3695__B _3693_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3751_ _3572_/Y _2984_/A _5321_/C _3750_/Y _3751_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_159_975 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4764__A2 _4757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_806 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2775__A1 _2735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_614 VGND VPWR sky130_fd_sc_hd__decap_12
X_2702_ _5357_/X _2690_/Y _2702_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_71_3 VGND VPWR sky130_fd_sc_hd__decap_6
X_3682_ _5522_/Q _3682_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_647 VGND VPWR sky130_fd_sc_hd__fill_2
X_5421_ _5421_/D data_out2[19] _4457_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_118_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_809 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_157 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_861 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_628 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_500 VGND VPWR sky130_fd_sc_hd__decap_12
X_5352_ _5351_/A _5351_/B _5352_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__4600__A _4600_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_200 VGND VPWR sky130_fd_sc_hd__fill_2
X_4303_ _4303_/A _4303_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_149 VGND VPWR sky130_fd_sc_hd__decap_4
X_5283_ _5252_/A _5252_/B _5515_/Q _5283_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5534__RESET_B _4322_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_929 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_417 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3216__A _3216_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_4234_ _4229_/X _4234_/B _4236_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_102_739 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_4165_ _4092_/X _4168_/B _4165_/C _4165_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_95_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_3116_ _3116_/A _3115_/X _3116_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_325 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2774__B _2774_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4096_ _4095_/X _4096_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_67_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_122 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5150__B _5149_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_807 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_667 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4047__A _5538_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3047_ _5463_/Q _3047_/B _3048_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_36_561 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3255__A2 _3253_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_712 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_199 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_380 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_918 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2790__A _2790_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_227 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_406 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4204__A1 data_in1[28] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3007__A2 _3004_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4998_ _4975_/X _4997_/X _4998_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_428 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3949_ _4664_/X _3950_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4755__A2 _4745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_945 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_444 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2803__A2_N _2802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_488 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4510__A _4504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_115 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_533 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5509__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5325__B _5325_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3126__A _4985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_130 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2965__A _2944_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_506 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4691__A1 _2733_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5341__A _4848_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3494__A2 _3480_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_303 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4691__B2 _4688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_678 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_83 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2693__B1_N _5351_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_829 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_43 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3246__A2 _3172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_892 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_339 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_745 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_87 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4994__A2 _4991_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_851 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_767 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_60 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_288 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_64 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_900 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2757__A1 _5300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_625 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5219__C _5218_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_282 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_945 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4123__C _4123_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_410 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_444 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_477 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4420__A _4422_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_487 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_894 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_498 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5171__A2 _4995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_447 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2859__B key_in[43] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_84 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5235__B key_in[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3036__A _2966_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_428 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4131__B1 _4718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4682__A1 _5514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4682__B2 _4677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_122 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_509 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5401__D _4797_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_615 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_881 VGND VPWR sky130_fd_sc_hd__decap_4
X_4921_ _4873_/A _4921_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_61_840 VGND VPWR sky130_fd_sc_hd__fill_2
X_4852_ _4852_/A _4851_/X _4852_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_61_884 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_361 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_737 VGND VPWR sky130_fd_sc_hd__fill_1
X_3803_ _3794_/Y _3802_/X _3794_/Y _3802_/X _3803_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_759 VGND VPWR sky130_fd_sc_hd__decap_4
X_4783_ _4043_/C _4781_/X data_out1[22] _4782_/X _5392_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_165_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_3734_ _3726_/Y _3733_/X _3734_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_119_625 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_3665_ _3661_/X _3728_/A _3665_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_617 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3533__A2_N _3532_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5404_ _4681_/X data_out2[2] _4477_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4330__A _4330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_680 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5162__A2 _5156_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2769__B _2767_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3596_ _3596_/A _3594_/X _3596_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_115_842 VGND VPWR sky130_fd_sc_hd__fill_2
X_5335_ _5334_/X _5309_/X _5335_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_38 VGND VPWR sky130_fd_sc_hd__fill_2
X_5266_ _5236_/A key_in[3] _5266_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4217_ _4215_/Y _4218_/B _4219_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_75_409 VGND VPWR sky130_fd_sc_hd__fill_2
X_5197_ _5197_/A _5252_/B _4679_/X _5197_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3476__A2 _3447_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_303 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_781 VGND VPWR sky130_fd_sc_hd__decap_3
X_4148_ _4100_/X _4132_/X _4107_/Y _4000_/Y _4131_/X _4149_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_141_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_859 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_280 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3881__C1 _3880_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_667 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_678 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_987 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_829 VGND VPWR sky130_fd_sc_hd__fill_1
X_4079_ _4077_/X _4078_/Y _4079_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3112__C _3037_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_380 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4976__A2 _4965_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2987__A1 _2984_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_0_0_clock_A clkbuf_4_1_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_158 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_46 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4505__A _4504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_715 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_68 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4189__B1 _4188_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_225 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_236 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_207 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_934 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3936__B1 _3935_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_720 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_411 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_282 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3400__A2 _3398_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_904 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_56 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5456__RESET_B _4415_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5336__A _5299_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_948 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5153__A2 _5147_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_958 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3164__A1 _4582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5481__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_396 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_193 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_258 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3058__A1_N _3128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2695__A _2695_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3467__A2 _3300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5071__A _5084_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_336 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_442 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3303__B _3303_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_902 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_892 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_391 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_542 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_147 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2978__A1 _2912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_169 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4415__A _4418_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_74 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_709 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4719__A2 _4712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4134__B _4106_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_770 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_741 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3973__B _3971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_797 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_628 VGND VPWR sky130_fd_sc_hd__decap_12
X_3450_ _3450_/A _3449_/Y _3450_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_171_745 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5144__A2 _5130_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_447 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_255 VGND VPWR sky130_fd_sc_hd__decap_12
X_3381_ _3342_/Y _3346_/Y _3341_/Y _3381_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_130_119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_5120_ _5121_/A _5119_/X _5122_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_111_300 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2902__A1 _4637_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_311 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2902__B2 _2901_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_344 VGND VPWR sky130_fd_sc_hd__fill_2
X_5051_ _5564_/Q _5038_/X _5051_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_878 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_770 VGND VPWR sky130_fd_sc_hd__fill_1
X_4002_ _3175_/Y _4001_/X _4002_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_37_100 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3213__B _3211_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_818 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_762 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_136 VGND VPWR sky130_fd_sc_hd__decap_12
X_4904_ _4914_/B _4902_/X _4904_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4325__A _4324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_501 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3091__B1 _3112_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_489 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_709 VGND VPWR sky130_fd_sc_hd__fill_2
X_4835_ _4802_/X _4842_/B _4834_/Y _4827_/A _4815_/X _4835_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_147_731 VGND VPWR sky130_fd_sc_hd__fill_1
X_4766_ _3870_/A _4757_/X data_out1[14] _4758_/X _4766_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_159_591 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3883__B _3878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_444 VGND VPWR sky130_fd_sc_hd__fill_1
X_3717_ _3788_/A _3715_/X _3716_/Y _3717_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_4697_ _2876_/A _4687_/X data_out2[11] _4688_/X _5413_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_20_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_734 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4060__A _4059_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3648_ _5290_/A _3646_/X _3647_/X _3651_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_136_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_778 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4995__A _4803_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_3579_ _3579_/A _3577_/X _3596_/A _3579_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_115_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_992 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_416 VGND VPWR sky130_fd_sc_hd__decap_12
X_5318_ _5317_/A _5317_/B _5319_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_88_534 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_491 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_867 VGND VPWR sky130_fd_sc_hd__decap_3
X_5249_ _5246_/X _5249_/B _5250_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_152_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_601 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_589 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3449__A2 _3410_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_697 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3404__A _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_100 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4219__B _4219_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3123__B _3122_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_902 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_689 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_979 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_467 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_311 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_312 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4235__A _4229_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_489 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_323 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_821 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_394 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3909__B1 _3908_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4889__B _4888_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3793__B _3776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_509 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_17 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_701 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5066__A _5037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_296 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3137__A1 _3074_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_469 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_255 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_288 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3688__A2 _3686_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4120__D _4119_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_512 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_81 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_910 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4924__A1_N _5554_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4129__B _4123_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_773 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3968__B _3945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2872__B _2822_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5377__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_456 VGND VPWR sky130_fd_sc_hd__fill_2
X_2950_ _2989_/A _2989_/B _2950_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_383 VGND VPWR sky130_fd_sc_hd__fill_2
X_2881_ _2852_/A _2879_/Y _2880_/X _2881_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_148_506 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5378__RESET_B _4507_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_876 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3984__A _3982_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4620_ _2707_/A _5301_/A VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5365__A2 _5363_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_742 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_904 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_550 VGND VPWR sky130_fd_sc_hd__fill_2
X_4551_ _5554_/Q _4547_/B _5554_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_144_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_937 VGND VPWR sky130_fd_sc_hd__decap_12
X_3502_ _3529_/A key_in[93] _3502_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4482_ _4477_/A _4482_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3208__B _3166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_918 VGND VPWR sky130_fd_sc_hd__decap_12
X_3433_ data_in2[26] _3391_/X _3393_/X _3432_/Y _5537_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_83_1010 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_320 VGND VPWR sky130_fd_sc_hd__fill_2
X_3364_ _3216_/A _3364_/B _4728_/X _3364_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_124_491 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_951 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_5103_ _5569_/Q _5102_/X _5569_/Q _5102_/X _5103_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4089__C1 _4088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3295_ _4639_/X _3291_/X _3292_/X _3293_/X _3294_/X _3295_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_98_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_921 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_686 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_5034_ _5034_/A _5031_/X _5034_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4039__B _4038_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_431 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_196 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3836__C1 _3835_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_423 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3878__B _3877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5053__B2 _5052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_264 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4055__A _4030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3597__C _3596_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_681 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2811__B1 _2783_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_342 VGND VPWR sky130_fd_sc_hd__decap_3
X_4818_ _5543_/Q _4837_/B _4818_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3367__A1 _3321_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_904 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_241 VGND VPWR sky130_fd_sc_hd__decap_3
X_4749_ _5327_/A _4745_/X data_out1[5] _4746_/X _5375_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_5_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_907 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4221__C _3368_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3118__B key_in[50] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_821 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_748 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_951 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_364 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_483 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_239 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_66 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2973__A _2973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_250 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4891__C _4890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_423 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_648 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_125 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3788__B _3786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_50 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_467 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_776 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_810 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_43 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_821 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_120 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_692 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_131 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5471__RESET_B _4396_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_142 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_803 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_153 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_898 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_313 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5400__RESET_B _4481_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_892 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_723 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3309__A _3287_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3028__B _3017_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_918 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_929 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_726 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_417 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4858__A1 _4848_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_450 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3044__A _2828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_312 VGND VPWR sky130_fd_sc_hd__decap_6
X_3080_ _4638_/X _3076_/X _3077_/X _3078_/X _3079_/X _3081_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_94_345 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3979__A _3966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2883__A _5355_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3294__B1 _3222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_968 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_294 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_754 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5559__RESET_B _4292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_456 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_979 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5035__A1 _4870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_916 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5035__B2 _4930_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_798 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3046__B1 _3042_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3982_ _3858_/Y _3981_/X _3982_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_22_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_949 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_804 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3210__C _3209_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2933_ _2934_/A key_in[13] _2933_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_15_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_837 VGND VPWR sky130_fd_sc_hd__decap_6
X_2864_ _2907_/A _2863_/X _2864_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4603__A _4605_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_4603_ _4605_/B _4603_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_163_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_701 VGND VPWR sky130_fd_sc_hd__decap_12
X_2795_ _4900_/A _2794_/B _2794_/X _2795_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_163_328 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3219__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4010__A2 _4008_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_892 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_4534_ _4533_/X _4542_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5137__C _5086_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4041__C _4041_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_233 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_862 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3760__B1_N _3759_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4465_ _4468_/A _4465_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_288 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_225 VGND VPWR sky130_fd_sc_hd__decap_8
X_3416_ _3416_/A _3415_/Y _3416_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3880__C _3879_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4396_ _4390_/X _4396_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3347_ _3342_/Y _3346_/Y _3342_/Y _3346_/Y _3347_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5542__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_995 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_634 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_38 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4992__B _4990_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3278_ _4720_/X _3274_/X _3354_/A _3284_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3889__A _3770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_5017_ _5017_/A _5017_/B _5017_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_250 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_924 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_710 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_220 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_47 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_776 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5026__B2 _5025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_253 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_415 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4785__B1 data_out1[23] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_24 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_982 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3713__B1_N _3693_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4513__A _4515_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_161 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_689 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_817 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4232__B _4214_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4001__A2 _5536_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3129__A _3129_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_704 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3760__A1 _3759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2968__A _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5344__A _5343_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_597 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3790__C _3804_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_640 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3512__A1 _3493_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_472 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_98 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3799__A _3797_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_721 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_42 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_916 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3311__B _3352_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_86 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_735 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4776__B1 data_out1[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_611 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4240__A2 _4227_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4423__A _4422_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_684 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5415__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_807 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_154 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4142__B _4142_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_520 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3200__B1 _3199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_553 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3751__A1 _3572_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2878__A _2878_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_501 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3751__B2 _3750_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5565__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5254__A _5243_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4172__A1_N _3287_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4250_ _4577_/A _4578_/A _4519_/X _4525_/X _4264_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_99_448 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_578 VGND VPWR sky130_fd_sc_hd__fill_2
X_3201_ _3188_/X _3200_/X _3188_/X _3200_/X _3201_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_802 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3503__A1 _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_109 VGND VPWR sky130_fd_sc_hd__decap_12
X_4181_ _4168_/Y _4182_/B _4183_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5404__D _4681_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3132_ _3107_/X _3163_/B _3107_/X _3163_/B _3133_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_868 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_367 VGND VPWR sky130_fd_sc_hd__decap_8
X_3063_ _3062_/A _3061_/X _3074_/A _3069_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_83_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_337 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3502__A _3529_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5393__RESET_B _4489_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_562 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_798 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_595 VGND VPWR sky130_fd_sc_hd__fill_2
X_3965_ _3954_/X _3964_/X _3954_/X _3964_/X _3965_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4333__A _4340_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2916_ _2998_/A _2916_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3896_ _3895_/A _3894_/X _3896_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5148__B _5148_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2793__A2 _2787_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2847_ _2847_/A _2847_/B _2847_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_148_166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3990__B2 _3989_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_2778_ _2778_/A _2777_/X _2778_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5566_ _5566_/D _5566_/Q _4284_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4987__B _4986_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3742__A1 _2717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_361 VGND VPWR sky130_fd_sc_hd__decap_8
X_4517_ _5436_/Q _4517_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_105_715 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2788__A _5301_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5497_ _5497_/D _5497_/Q _4366_/X _5429_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5164__A _5478_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_759 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_556 VGND VPWR sky130_fd_sc_hd__decap_3
X_4448_ _4469_/A _4449_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_59 VGND VPWR sky130_fd_sc_hd__decap_12
X_4379_ _4381_/A _4379_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_59_824 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_781 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_492 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_431 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5247__A1 _4679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_879 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4508__A _4504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2954__C _2953_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_36 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3412__A _5472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_68 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_231 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_916 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3131__B _3131_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_938 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_34 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5438__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_34 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2970__B key_in[78] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4222__A2 _4211_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_943 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3964__A1_N _3131_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4243__A _4241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_965 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_790 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_453 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3981__A1 _3770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3981__B2 _3980_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_614 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_520 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_647 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_629 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2698__A _5252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_168 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_821 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_718 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_898 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_589 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_886 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3497__B1 _3466_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_665 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5238__A1 _4636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5238__B2 _5237_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_613 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4418__A _4418_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_326 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3322__A _3322_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_754 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_540 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_253 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_562 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3041__B key_in[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_713 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_893 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_532 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_757 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4749__B1 data_out1[5] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2880__B _2921_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5249__A _5246_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3750_ _5525_/Q _3750_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_289 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3695__C _3694_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3421__B1 _3436_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_442 VGND VPWR sky130_fd_sc_hd__fill_2
X_2701_ _3603_/B _2723_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2775__A2 _2774_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_3681_ _3681_/A _3680_/X _3681_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_146_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_103 VGND VPWR sky130_fd_sc_hd__decap_12
X_5420_ _5420_/D data_out2[18] _4458_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_64_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_851 VGND VPWR sky130_fd_sc_hd__decap_3
X_5351_ _5351_/A _5351_/B _5351_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_372 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4600__B _4600_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_512 VGND VPWR sky130_fd_sc_hd__decap_6
X_4302_ _4303_/A _4302_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_320 VGND VPWR sky130_fd_sc_hd__fill_2
X_5282_ data_in2[3] _5222_/X _5252_/X _5281_/X _5514_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_141_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_876 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_4233_ _4230_/X _4233_/B _4232_/Y _4234_/B VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_59_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3216__B _3143_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_217 VGND VPWR sky130_fd_sc_hd__decap_8
X_4164_ _4158_/X _4163_/B _4165_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_68_654 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5574__RESET_B _4273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_440 VGND VPWR sky130_fd_sc_hd__decap_8
X_3115_ _3112_/X _3115_/B _3115_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_68_698 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4328__A _4330_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4095_ _4094_/X _4095_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5503__RESET_B _4358_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_134 VGND VPWR sky130_fd_sc_hd__decap_4
X_3046_ _4637_/X _3040_/X _3041_/X _3042_/X _3045_/X _3047_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_82_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_551 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_882 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_0_0_clock_A clkbuf_2_0_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_718 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_392 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_543 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2790__B key_in[73] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_565 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4204__A2 _4125_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4997_ _4555_/A _4965_/X _4997_/C _4987_/A _4997_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_23_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5159__A _5159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4063__A _4014_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_442 VGND VPWR sky130_fd_sc_hd__decap_12
X_3948_ data_in1[17] _3837_/X _3929_/X _3947_/Y _5496_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_139_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4998__A _4975_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3879_ _3873_/Y _3877_/X _3879_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_164_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_862 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_617 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_5549_ _4545_/X _4545_/A _4303_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3407__A _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_353 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3126__B _3081_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_632 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_548 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_963 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_142 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2965__B _2965_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_762 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4691__A2 _4687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5341__B _5341_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_808 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_540 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4979__B1 _4978_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_860 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_882 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2981__A _2998_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__A3 _4992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_841 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5069__A _5068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_32 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2757__A2 key_in[104] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_76 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_985 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_957 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4701__A _4701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5156__B1 _4573_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_456 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_692 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3317__A _2885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3036__B _3036_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_898 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_695 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_91 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4131__A1 _3905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_559 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4131__B2 _3520_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_451 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4682__A2 _4674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2693__A1 _5321_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_849 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3052__A _3052_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_540 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_627 VGND VPWR sky130_fd_sc_hd__decap_12
X_4920_ _2907_/A _4925_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2891__A _2714_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_852 VGND VPWR sky130_fd_sc_hd__fill_2
X_4851_ _5548_/Q _4850_/X _5548_/Q _4850_/X _4851_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_896 VGND VPWR sky130_fd_sc_hd__decap_12
X_3802_ _3795_/X _3801_/X _3802_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_20_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_4782_ _4700_/A _4782_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_248 VGND VPWR sky130_fd_sc_hd__fill_2
X_3733_ _3705_/Y _3727_/Y _3731_/X _3732_/Y _3733_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_146_423 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4611__A _4610_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3664_ _3663_/X _3728_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_5403_ _5403_/D data_out2[1] _4478_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_415 VGND VPWR sky130_fd_sc_hd__fill_2
X_3595_ _3596_/A _3594_/X _3595_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_821 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2769__C _5310_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3227__A _3227_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5334_ _4836_/A _5334_/B _5334_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_170_982 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_204 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_515 VGND VPWR sky130_fd_sc_hd__decap_4
X_5265_ _5234_/A key_in[35] _5265_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_141_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_857 VGND VPWR sky130_fd_sc_hd__fill_2
X_4216_ _4231_/A _4203_/B _4218_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_259 VGND VPWR sky130_fd_sc_hd__fill_2
X_5196_ data_in2[0] _4574_/B _5175_/X _5195_/X _5196_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_18_15 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3330__C1 _3329_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_315 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_933 VGND VPWR sky130_fd_sc_hd__decap_12
X_4147_ _3395_/X _4145_/X _4146_/X _4147_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_55_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3881__B1 _3857_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_646 VGND VPWR sky130_fd_sc_hd__fill_1
X_4078_ _3955_/Y _4076_/X _4078_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3897__A _3895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_318 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_627 VGND VPWR sky130_fd_sc_hd__fill_2
X_3029_ _2999_/A _3028_/X _3060_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_392 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2987__A2 _2984_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4189__A1 _3316_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3936__A1 _3075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_4_0_clock_A clkbuf_4_5_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_219 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_103 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_793 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4521__A _4521_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_24 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_979 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_147 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_776 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_478 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5336__B key_in[37] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_68 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_117 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_990 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5153__A3 _5140_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_436 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_459 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3164__A2 _3163_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_960 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5496__RESET_B _4367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_705 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_876 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5018__B1_N _5017_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2976__A _4943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_226 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5425__RESET_B _4452_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5352__A _5351_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_345 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_879 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2695__B _2695_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5071__B _5085_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_771 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_21 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_83 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5502__D _4089_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_104 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_510 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_690 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3600__A _3600_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_31 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_863 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2978__A2 _2975_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_682 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_598 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_209 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_557 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_935 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_581 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_957 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4431__A _4426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_905 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_786 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3047__A _5463_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_3380_ _5472_/Q _3379_/B _3413_/B _3414_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_170_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_970 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2902__A2 _2898_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_470 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2886__A _5523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3165__A1_N _3162_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_226 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5262__A _3626_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5050_ _5037_/X _5052_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_579 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_4001_ _3062_/A _5536_/Q _5527_/Q _4000_/Y _4001_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_66_933 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5412__D _4695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_646 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_281 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_432 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_657 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_785 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_318 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4606__A _4605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3510__A _3510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_148 VGND VPWR sky130_fd_sc_hd__decap_4
X_4903_ _4914_/B _4902_/X _4903_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_33_351 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3091__B2 _3090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_513 VGND VPWR sky130_fd_sc_hd__decap_4
X_4834_ _4833_/A _4833_/B _4834_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_21_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_507 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_721 VGND VPWR sky130_fd_sc_hd__fill_2
X_4765_ _2797_/A _3870_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4341__A _4341_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_905 VGND VPWR sky130_fd_sc_hd__decap_8
X_3716_ _3712_/X _3714_/Y _3716_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4696_ _5522_/Q _2876_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_135_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_264 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_489 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_949 VGND VPWR sky130_fd_sc_hd__fill_2
X_3647_ _5290_/A _3646_/X _3647_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_106_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_746 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_128 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_49 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_139 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_960 VGND VPWR sky130_fd_sc_hd__fill_2
X_3578_ _3578_/A _3575_/X _3596_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_513 VGND VPWR sky130_fd_sc_hd__decap_6
X_5317_ _5317_/A _5317_/B _5319_/B VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_103_824 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_428 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5172__A _5172_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_5248_ _5246_/X _5249_/B _5278_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_152_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_47 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3404__B key_in[58] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_410 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_944 VGND VPWR sky130_fd_sc_hd__fill_2
X_5179_ _3577_/A _3578_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4219__C _4218_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_966 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_958 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4516__A _4515_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3606__B1 _3619_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_852 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_302 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4235__B _4234_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_479 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3082__A1 _4985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_324 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_41 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_335 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_507 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_85 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_529 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3909__A1 _3062_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_528 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4251__A _4517_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5066__B _5065_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_723 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3594__A2_N _3593_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3137__A2 _3096_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_971 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_789 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_161 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_288 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5082__A _5081_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_579 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4098__B1 _3175_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_922 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_687 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_101 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_97 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3845__B1 _3817_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4426__A _4419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_830 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3968__C _3924_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_874 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_479 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_822 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_833 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2820__A1 _2819_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2880_ _2855_/Y _2921_/B _2880_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_181 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_332 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3984__B _3983_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_899 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5257__A _2716_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_398 VGND VPWR sky130_fd_sc_hd__decap_4
X_4550_ _5553_/Q _4541_/B _5553_/D VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_562 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_253 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_798 VGND VPWR sky130_fd_sc_hd__fill_1
X_3501_ _3501_/A key_in[29] _3501_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_949 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5407__D _5407_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4481_ _4477_/A _4481_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_3432_ _3317_/X _3432_/B _3432_/C _3432_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_143_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_310 VGND VPWR sky130_fd_sc_hd__fill_1
X_3363_ data_in2[24] _3172_/X _3316_/X _3362_/Y _3363_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_112_621 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_866 VGND VPWR sky130_fd_sc_hd__decap_3
X_5102_ _5037_/X _5101_/X _5102_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_140_963 VGND VPWR sky130_fd_sc_hd__decap_12
X_3294_ _3291_/A key_in[119] _3222_/X _3294_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_58_719 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4089__B1 _4071_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_527 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_933 VGND VPWR sky130_fd_sc_hd__fill_2
X_5033_ _5030_/Y _5032_/Y _5033_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3836__B1 _3812_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_616 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4336__A _4339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_619 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_800 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4055__B _4053_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_49 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5053__A2_N _5052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_693 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2811__A1 data_in2[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5471__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_866 VGND VPWR sky130_fd_sc_hd__decap_12
X_4817_ _4817_/A _4821_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_166_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5167__A _5167_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_220 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4071__A _4026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3367__A2 _3349_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4748_ _5181_/B _5327_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_275 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_4679_ _3588_/A _4679_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_418 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_429 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_737 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_941 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3415__A _3412_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_866 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1000 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3827__B1 _3826_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_903 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2973__B _2972_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_262 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4246__A _4246_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3788__C _3787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_744 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3958__B1_N _3957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_118 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_129 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_121 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_66 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_143 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_154 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_849 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_877 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_176 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5077__A _5566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_359 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3309__B _3309_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_735 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5440__RESET_B _4434_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4858__A2 _4847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_598 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_226 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3325__A _3324_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5131__A1_N _5571_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_462 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_218 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_91 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3979__B _3972_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3294__A1 _3291_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4156__A _4155_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3060__A _3060_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5494__CLK _5430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5035__A2 _5033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_232 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_541 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_608 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3046__A1 _4637_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3046__B2 _3045_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3981_ _3770_/Y _5535_/Q _3020_/A _3980_/Y _3981_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3995__A _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_2932_ _2968_/A key_in[45] _2932_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_94_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_326 VGND VPWR sky130_fd_sc_hd__decap_8
X_2863_ _4637_/X _2859_/X _2860_/X _2861_/X _2862_/X _2863_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_148_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5528__RESET_B _4329_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_696 VGND VPWR sky130_fd_sc_hd__decap_12
X_4602_ _4602_/A _4605_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_129_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_2794_ _5456_/Q _2794_/B _2794_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_7_50 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_713 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3219__B key_in[21] VGND VPWR sky130_fd_sc_hd__diode_2
X_4533_ _4529_/X _4533_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_757 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_391 VGND VPWR sky130_fd_sc_hd__decap_8
X_4464_ _4468_/A _4464_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_429 VGND VPWR sky130_fd_sc_hd__decap_12
X_3415_ _3412_/X _3413_/X _3414_/Y _3415_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_4395_ _4390_/X _4395_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3235__A _3233_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3346_ _3343_/X _3344_/X _3345_/Y _3346_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_113_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_869 VGND VPWR sky130_fd_sc_hd__decap_4
X_3277_ _3288_/A _3354_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3439__A2_N _4791_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3889__B _3887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_903 VGND VPWR sky130_fd_sc_hd__fill_2
X_5016_ _5562_/Q _5015_/X _5562_/Q _5015_/X _5017_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_26_402 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_788 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_265 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_107 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4785__A1 _4784_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4785__B2 _4782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2796__B1 _2785_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_47 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_348 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4232__C _4232_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_189 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3129__B _3127_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_724 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_234 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3760__A2 _3758_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2968__B key_in[46] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3145__A _3043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3512__A2 _3539_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_985 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2720__B1 _2744_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_484 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2984__A _2984_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_357 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3799__B _3799_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_733 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5510__D _4249_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_744 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_906 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_54 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_777 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_980 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_747 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4776__A1 _4775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4776__B2 _4770_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_641 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_623 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_696 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_122 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_184 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4142__C _4142_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_381 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3200__A1 _3199_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_851 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3751__A2 _2984_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_862 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_405 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2878__B _2920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_204 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2773__A1_N _2736_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4154__A2_N _4153_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3055__A _2910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3200_ _3199_/A _3198_/Y _3199_/Y _3200_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3503__A2 key_in[125] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_760 VGND VPWR sky130_fd_sc_hd__decap_3
X_4180_ _4178_/X _4196_/B _4182_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_814 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_622 VGND VPWR sky130_fd_sc_hd__decap_12
X_3131_ _3131_/A _3131_/B _3163_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__2894__A _2822_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5270__A _4827_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3062_ _3062_/A _3061_/X _3074_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_94_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_305 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_711 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3502__B key_in[93] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_593 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5420__D _5420_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0_0_clock_A clkbuf_2_1_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_872 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_788 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_416 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_894 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_991 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4614__A _4525_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3964_ _3131_/B _3963_/X _3131_/B _3963_/X _3964_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3975__C1 _3974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2915_ _2915_/A _2914_/X _2998_/A VGND VPWR sky130_fd_sc_hd__xor2_4
X_3895_ _3895_/A _3894_/X _3895_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_148_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_808 VGND VPWR sky130_fd_sc_hd__fill_2
X_2846_ _2778_/X _2846_/B _2849_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2793__A3 _2789_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_189 VGND VPWR sky130_fd_sc_hd__fill_2
X_5565_ _4564_/X _5065_/A _4285_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2777_ _2723_/A _2723_/B _2776_/X _2777_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_145_841 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_554 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3742__A2 _3710_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4516_ _4515_/A _4516_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5496_ _5496_/D _2889_/A _4367_/X _5429_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1004 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_738 VGND VPWR sky130_fd_sc_hd__fill_2
X_4447_ _4267_/Y _4469_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_803 VGND VPWR sky130_fd_sc_hd__decap_3
X_4378_ _4381_/A _4378_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_313 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_3329_ _3259_/A _3304_/X _3258_/Y _3329_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_112_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_346 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5180__A _5327_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_443 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5247__A2 _5215_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_176 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3412__B _3379_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_850 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_202 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_427 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_449 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4524__A _4524_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_421 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_983 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4243__B _4242_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4862__A1_N _4545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3981__A2 _5535_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3718__C1 _3717_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_626 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5355__A _5355_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3194__B1 _5023_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2698__B _2698_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_61 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2941__B1 _3759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_855 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5505__D _4166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4143__C1 _4142_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_888 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_760 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3497__A1 _3155_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3497__B2 _3468_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_493 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5090__A _5472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3603__A _3603_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_806 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_143 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5238__A2 _5234_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_809 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_232 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_168 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_596 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4749__A1 _5327_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4749__B2 _4746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4434__A _4438_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_769 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5249__B _5249_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_955 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3421__B2 _3420_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5532__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_791 VGND VPWR sky130_fd_sc_hd__fill_2
X_2700_ _5518_/Q _3603_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3680_ _3680_/A _3669_/X _3680_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_115 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2889__A _2889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5265__A _5234_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5350_ _5350_/A _5319_/C _5351_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_57_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4301_ _4303_/A _4301_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_5281_ _5281_/A _5281_/B _5281_/C _5281_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5415__D _5415_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_192 VGND VPWR sky130_fd_sc_hd__decap_12
X_4232_ _4195_/X _4214_/X _4232_/C _4232_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3216__C _4718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4685__B1 data_out2[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_942 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4609__A _4646_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4163_ _4158_/X _4163_/B _4168_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3513__A _3513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_752 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_677 VGND VPWR sky130_fd_sc_hd__fill_2
X_3114_ _3033_/Y _3088_/X _3113_/X _3115_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_95_463 VGND VPWR sky130_fd_sc_hd__fill_2
X_4094_ _4073_/X _4093_/X _4094_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_647 VGND VPWR sky130_fd_sc_hd__fill_2
X_3045_ _3043_/X key_in[112] _3044_/X _3045_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_167_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_894 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5543__RESET_B _4310_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_202 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_213 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4344__A _4341_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4996_ _4996_/A _5000_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_23_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5159__B _5159_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_419 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3948__C1 _3947_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4063__B _4038_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_clock_A clkbuf_2_2_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3947_ _3835_/A _3945_/Y _3947_/C _3947_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_51_599 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_454 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_49 VGND VPWR sky130_fd_sc_hd__decap_12
X_3878_ _3873_/Y _3877_/X _3878_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4998__B _4997_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_975 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_498 VGND VPWR sky130_fd_sc_hd__fill_2
X_2829_ _2859_/A key_in[106] _2828_/X _2829_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__2799__A _2799_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5175__A _5197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4912__A1 _4911_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5548_ _5548_/D _5548_/Q _4305_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_155_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_896 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_490 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_395 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_5479_ _3580_/X _3577_/A _4387_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_644 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4519__A _4518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_430 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_741 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_806 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2965__C _2964_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3423__A _3422_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_68 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5405__CLK _5402_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_463 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_316 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3240__A2_N _3239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_198 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_284 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4979__A1 _4974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_530 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_850 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2981__B _2998_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_680 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5555__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_207 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_864 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_11 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_73 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__A1 _3400_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_739 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_780 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_796 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_88 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_947 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_115 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_969 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_71 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_434 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5156__B2 _5155_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5085__A _5072_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_660 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_800 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_31 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_885 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_192 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1009 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_354 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3823__A2_N _3822_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3036__C _2965_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_516 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_227 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4131__A2 _5541_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4429__A _4426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_901 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2693__A2 _5348_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_338 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3052__B _3052_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_308 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2891__B _2891_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_831 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_533 VGND VPWR sky130_fd_sc_hd__fill_2
X_4850_ _4819_/A _4849_/X _4850_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_127_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4164__A _4158_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_555 VGND VPWR sky130_fd_sc_hd__fill_2
X_3801_ _3801_/A _3820_/B _3801_/X VGND VPWR sky130_fd_sc_hd__xor2_4
X_4781_ _4672_/X _4781_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_14_780 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_774 VGND VPWR sky130_fd_sc_hd__fill_2
X_3732_ _3661_/X _3730_/A _3642_/X _3732_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_119_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_785 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5147__A1 _5143_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3663_ _3662_/X _3663_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_5402_ _5402_/D data_out2[0] _4479_/X _5402_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3594_ _3583_/C _3593_/X _3583_/C _3593_/X _3594_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_129 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3227__B _3226_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5333_ _5325_/X _5332_/X _5325_/X _5332_/X _5333_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_717 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5428__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_5264_ _4817_/A _5238_/X _5241_/X _5264_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_141_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_4215_ _4214_/X _4215_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_4_11_0_clock_A clkbuf_3_5_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_549 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4339__A _4339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_441 VGND VPWR sky130_fd_sc_hd__fill_1
X_5195_ _5281_/A _5192_/X _5194_/X _5195_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3243__A _3244_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3330__B1 _3304_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_463 VGND VPWR sky130_fd_sc_hd__decap_12
X_4146_ _3394_/Y _4145_/X _4146_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_411 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3881__A1 data_in1[14] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_49 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5578__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_455 VGND VPWR sky130_fd_sc_hd__fill_2
X_4077_ _3955_/Y _4076_/X _4077_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3348__A1_N _3333_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5083__B1 _5082_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3897__B _3896_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3028_ _2999_/B _3017_/X _3028_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_70_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_505 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_544 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4074__A _4045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_853 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_205 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4189__A2 _5539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4979_ _4974_/Y _4978_/B _4978_/Y _4982_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4802__A _4857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3936__A2 _3933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_947 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_115 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_446 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3149__B1 _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_916 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_clock_A clkbuf_4_9_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_800 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_298 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_844 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_630 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_641 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_332 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2976__B _2936_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_696 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5352__B _5351_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_357 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_560 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_625 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5465__RESET_B _4403_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_95 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2992__A _3065_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5074__B1 _5073_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_308 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3194__A2_N _3228_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_522 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3600__B _3592_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_43 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_560 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_700 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4712__A _4699_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_424 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5110__B1_N _5109_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_221 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_969 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_446 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_917 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3328__A _3304_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_405 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_660 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_107 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3132__A2_N _3163_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4888__B1 _4875_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_80 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3047__B _3047_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3560__B1 _4791_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_674 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2902__A3 _2899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_825 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_493 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5262__B _5262_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_335 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4159__A _4112_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4000_ _5536_/Q _4000_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_614 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3777__A2_N _3776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_411 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3998__A _3903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_168 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_105 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3510__B _3510_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4902_ _4885_/Y _4889_/Y _4902_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_4833_ _4833_/A _4833_/B _4842_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_525 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4622__A _2934_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4764_ _3875_/A _4757_/X data_out1[13] _4758_/X _4764_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_147_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_3715_ _3712_/X _3714_/Y _3715_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4695_ _2842_/A _4687_/X data_out2[10] _4688_/X _4695_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_101_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_3646_ _3635_/Y _3645_/X _3635_/Y _3645_/X _3646_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_630 VGND VPWR sky130_fd_sc_hd__decap_12
X_3577_ _3577_/A _3600_/A _3577_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_652 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3272__A1_N _3268_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5316_ _5276_/X _5281_/B _5317_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_142_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_15 VGND VPWR sky130_fd_sc_hd__decap_8
X_5247_ _4679_/X _5215_/X _5217_/X _5249_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XANTENNA__4069__A _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_666 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_5178_ _3573_/A _5178_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_29_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1018 VGND VPWR sky130_fd_sc_hd__fill_2
X_4129_ _4128_/X _4123_/B _4129_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_29_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_809 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3701__A _3680_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_488 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3606__B2 _3605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_149 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_864 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_190 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_303 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_650 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3082__A2 _3081_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_314 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_324 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_325 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_335 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_336 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3909__A2 _3906_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_530 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4251__B _4668_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2939__A2_N _2938_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3148__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_758 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_408 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_50 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_983 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_536 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5513__D _5513_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4098__A1 _3175_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4098__B2 _4097_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_974 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3845__A1 _3818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_411 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_891 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_956 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4707__A _4707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_455 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3611__A _3609_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_680 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_778 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2820__A2 _2819_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_193 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4442__A _4443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_733 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_210 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_540 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3500_ _3528_/A key_in[61] _3500_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_156_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_562 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3781__B1 _3828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_725 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_4480_ _4477_/A _4480_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_747 VGND VPWR sky130_fd_sc_hd__decap_4
X_3431_ _3431_/A _3431_/B _3432_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_143_257 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_801 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3533__B1 _5154_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_3362_ _3317_/X _3362_/B _3362_/C _3362_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__5387__RESET_B _4496_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5101_ _5568_/Q _5091_/X _5101_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_3_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_333 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_975 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4089__A1 data_in1[23] VGND VPWR sky130_fd_sc_hd__diode_2
X_3293_ _3293_/A key_in[87] _3293_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5423__D _4719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_5032_ _5031_/X _5032_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3836__A1 data_in1[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_967 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_230 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_764 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4617__A _5203_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_550 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3521__A _3520_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_499 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_594 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_691 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_469 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4055__C _4054_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_119 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_834 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2811__A2 _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_480 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_193 VGND VPWR sky130_fd_sc_hd__decap_12
X_4816_ _4802_/X _4823_/B _4814_/Y _5448_/Q _4815_/X _4816_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4352__A _4349_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_878 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_355 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5210__B1 _4811_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5167__B _5167_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4747_ _5287_/A _4745_/X data_out1[4] _4746_/X _5374_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4071__B _3950_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_27 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_49 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3669__A2_N _3668_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4678_ _3573_/A _4674_/X data_out2[0] _4677_/X _5402_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_162_544 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_3629_ _3630_/A _3628_/X _3631_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5183__A _5203_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3524__B1 _3396_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_26 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_845 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_493 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3415__B _3413_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_709 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_400 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1012 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_496 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3827__A1 _2714_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_591 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4841__B1_N _4840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_753 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3607__A2_N _3606_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4527__A _4577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_509 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5029__B1 _5028_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3431__A _3431_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_116 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4246__B _4246_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_756 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4226__B1_N _4225_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_981 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_299 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5358__A _5358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_155 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_867 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_816 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_316 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_827 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4262__A _4631_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_327 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_177 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5201__B1 _3583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_188 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_199 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5077__B _5065_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_552 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5508__D _5508_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_408 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5480__RESET_B _4386_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_815 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5268__B1 _5303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_474 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_848 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3818__A1 _2918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4437__A _4438_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3341__A _3340_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3294__A2 key_in[119] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_403 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_1_0_0_clock_A clkbuf_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_745 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3060__B _3060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5035__A3 _5034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_553 VGND VPWR sky130_fd_sc_hd__decap_12
X_3980_ _5535_/Q _3980_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3046__A2 _3040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3995__B _3993_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_597 VGND VPWR sky130_fd_sc_hd__decap_12
X_2931_ _2905_/Y _2913_/X _2931_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_16_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_299 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_817 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_130 VGND VPWR sky130_fd_sc_hd__fill_1
X_2862_ _2859_/A key_in[107] _2828_/X _2862_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_87_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_349 VGND VPWR sky130_fd_sc_hd__decap_8
X_4601_ _5443_/Q _4601_/B _4602_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__5418__D _4709_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2793_ _4637_/A _2787_/X _2789_/X _2790_/X _2792_/X _2794_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_144_500 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_574 VGND VPWR sky130_fd_sc_hd__decap_12
X_4532_ _4517_/Y _4531_/X mode _4531_/X _4532_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_156_371 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4900__A _4900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_831 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5568__RESET_B _4281_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_95 VGND VPWR sky130_fd_sc_hd__fill_2
X_4463_ _4468_/A _4463_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3516__A _3516_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3414_ _3342_/Y _3414_/B _3346_/Y _3414_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_144_599 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_920 VGND VPWR sky130_fd_sc_hd__fill_2
X_4394_ _4390_/X _4394_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_931 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3235__B _3258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_430 VGND VPWR sky130_fd_sc_hd__decap_12
X_3345_ _3268_/Y _3297_/X _3271_/X _3345_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__5259__B1 _5230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_772 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_837 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_614 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_474 VGND VPWR sky130_fd_sc_hd__fill_2
X_3276_ _3275_/X _3288_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_5015_ _4975_/X _5014_/X _5015_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_73_509 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4347__A _4340_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3251__A _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_786 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_937 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_414 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4967__A2_N _4966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_959 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_918 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3593__A2_N _3592_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_575 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_277 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_981 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_992 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4785__A2 _4781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5178__A _3573_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_642 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2796__B2 _2795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_647 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_848 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_59 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_861 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4810__A _4837_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3129__C _3128_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_736 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_842 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_875 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3426__A _3361_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_953 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_141 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4150__B1_N _4173_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_975 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2720__B2 _2719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_794 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2984__B _2984_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_369 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_892 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_531 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_255 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4776__A2 _4769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_759 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3433__C1 _3432_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5088__A _5087_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_951 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_664 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_657 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_9 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3736__B1 _3735_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4720__A _4720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3200__A2 _3198_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_149 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3336__A _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3055__B _3055_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4161__B1 _4138_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_314 VGND VPWR sky130_fd_sc_hd__decap_12
X_3130_ _3125_/Y _3129_/Y _3125_/Y _3129_/Y _3131_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5461__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_634 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2894__B _2871_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_945 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5270__B _5270_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_590 VGND VPWR sky130_fd_sc_hd__decap_12
X_3061_ _3060_/A _3060_/B _3060_/X _3061_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__4167__A _4126_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_689 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3071__A _2927_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_723 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_211 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5067__A2_N _5066_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_756 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_981 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_225 VGND VPWR sky130_fd_sc_hd__decap_4
X_3963_ _3958_/X _3962_/X _3963_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__4614__B _4629_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_603 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_247 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3975__B1 _3950_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2914_ _2913_/A _2912_/X _2913_/X _2914_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_149_636 VGND VPWR sky130_fd_sc_hd__fill_2
X_3894_ _3885_/Y _3893_/X _3885_/Y _3893_/X _3894_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_2845_ _2842_/A _2842_/B _2844_/Y _2850_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_164_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_116 VGND VPWR sky130_fd_sc_hd__decap_6
X_5564_ _4563_/X _5564_/Q _4286_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4630__A _4630_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2776_ _2776_/A _2726_/A _2776_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_853 VGND VPWR sky130_fd_sc_hd__fill_1
X_4515_ _4515_/A _4515_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5495_ _3928_/X _3902_/C _4368_/X _5429_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_503 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3009__A1_N _3050_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_683 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1016 VGND VPWR sky130_fd_sc_hd__decap_4
X_4446_ _4443_/A _4446_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_962 VGND VPWR sky130_fd_sc_hd__fill_2
X_4377_ _4381_/A _4377_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_601 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_3328_ _3304_/A _3328_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_422 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_37 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_550 VGND VPWR sky130_fd_sc_hd__decap_6
X_3259_ _3259_/A _3258_/Y _3305_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_74_829 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4077__A _3955_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_520 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_862 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_778 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4805__A _4805_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_350 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_715 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_47 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_912 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_400 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_258 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_601 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_483 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5419__RESET_B _4459_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_105 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3718__B1 _3699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4540__A _4837_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_864 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3194__B2 _3228_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_875 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_672 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2698__C _5518_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_886 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4229__A2_N _4228_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5145__A1_N _4572_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_683 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2941__A1 _2799_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_525 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2941__B2 _3110_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5484__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_599 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_558 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4143__B1 _4127_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3497__A2 _3466_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_99 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_591 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3603__B _3603_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_21 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5238__A3 _5235_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5521__D _2853_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_60 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4715__A _5530_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_277 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4749__A2 _4745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_247 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_556 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_781 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_989 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3709__B1 _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_476 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4450__A _4449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_487 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5265__B key_in[35] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_864 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_801 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3066__A _2991_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4300_ _4303_/A _4300_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_127_897 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_660 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_171 VGND VPWR sky130_fd_sc_hd__fill_2
X_5280_ _5277_/X _5280_/B _5281_/C VGND VPWR sky130_fd_sc_hd__nand2_4
X_4231_ _4231_/A _4213_/X _4233_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_4_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4685__A1 _5321_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5281__A _5281_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_74 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4685__B2 _4677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4999__A1_N _4559_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_399 VGND VPWR sky130_fd_sc_hd__decap_12
X_4162_ _4159_/X _4198_/A _4163_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4609__B _4609_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3113_ _3113_/A _3088_/B _3113_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_4093_ _4074_/X _4082_/X _4093_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_306 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5431__D _5431_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_339 VGND VPWR sky130_fd_sc_hd__decap_12
X_3044_ _2828_/X _3044_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_309 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4625__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_191 VGND VPWR sky130_fd_sc_hd__decap_12
X_4995_ _4803_/Y _4995_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_51_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_269 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3948__B1 _3929_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4070__C1 _4069_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3946_ _3945_/A _3945_/B _3947_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3563__A1_N _3557_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_466 VGND VPWR sky130_fd_sc_hd__decap_12
X_3877_ _3874_/X _3876_/Y _3877_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__5512__RESET_B _4348_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_937 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4360__A _4354_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2828_ _2828_/A _2828_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2799__B _2799_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5175__B _5252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_853 VGND VPWR sky130_fd_sc_hd__decap_3
X_5547_ _5547_/D _5547_/Q _4306_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2759_ _4882_/A _2759_/B _2759_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4912__A2 _4910_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_300 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_525 VGND VPWR sky130_fd_sc_hd__decap_6
X_5478_ _5171_/X _5478_/Q _4388_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_867 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_878 VGND VPWR sky130_fd_sc_hd__decap_12
X_4429_ _4426_/X _4429_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_770 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3704__A _3603_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2687__B1 _2686_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_943 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_188 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4979__A2 _4978_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4535__A _5543_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_704 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_169 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_692 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_180 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2772__A1_N _2753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_219 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_52 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_876 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__A2 _3401_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_85 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_230 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_792 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_617 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_291 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_403 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5366__A _5299_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_274 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4270__A _4271_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_127 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_842 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3167__A1 _3143_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_446 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5085__B _5085_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5516__D _5354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_992 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2914__A1 _2913_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_897 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_480 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_924 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_935 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_497 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_467 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_564 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4445__A _4443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_895 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_692 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4164__B _4163_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_865 VGND VPWR sky130_fd_sc_hd__fill_2
X_3800_ _3799_/X _3820_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_4780_ _3085_/A _4043_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_159_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_770 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_792 VGND VPWR sky130_fd_sc_hd__decap_12
X_3731_ _3666_/A _3661_/X _3730_/Y _3731_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_9_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5276__A _5253_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4180__A _4178_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_959 VGND VPWR sky130_fd_sc_hd__decap_3
X_3662_ _5516_/Q _3659_/X _3662_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5147__A2 _5145_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_149 VGND VPWR sky130_fd_sc_hd__decap_4
X_5401_ _4797_/X data_out1[31] _4480_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_406 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5426__D _5426_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3593_ _3587_/X _3592_/Y _3587_/X _3592_/Y _3593_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_812 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5332_ _5332_/A _5332_/B _5332_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_480 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_5263_ _5260_/A _5261_/A _5262_/X _5263_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_125_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_4214_ _4794_/X _4212_/X _4213_/X _4214_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_141_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_420 VGND VPWR sky130_fd_sc_hd__decap_12
X_5194_ _3573_/A _5226_/A _5194_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3330__A1 _3254_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_762 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3243__B _3244_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4145_ _3932_/Y _5542_/Q _4720_/X _3548_/Y _4145_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_84_924 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_475 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3881__A2 _3837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_328 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_clock_A clkbuf_3_7_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4076_ _3858_/Y _5539_/Q _3143_/C _3463_/Y _4076_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_95_294 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_136 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5083__A1 _5076_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_478 VGND VPWR sky130_fd_sc_hd__fill_2
X_3027_ _5527_/Q _3062_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3094__B1 _3176_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4355__A _4354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2841__B1 _2815_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4074__B _4057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_556 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_364 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_217 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4978_ _4974_/Y _4978_/B _4978_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_11_228 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_915 VGND VPWR sky130_fd_sc_hd__fill_2
X_3929_ _3839_/A _3812_/B _3113_/A _3929_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_137_403 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5186__A _4635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4090__A _4664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_458 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3149__A1 _3145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_469 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_928 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_620 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_834 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_24 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_377 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3434__A _3519_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_388 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4829__A1_N _4542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_369 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5522__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_550 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_924 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_784 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3773__B1_N _3819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_946 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_434 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2992__B _2991_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_445 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_968 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5074__A1 _5071_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_383 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_534 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5434__RESET_B _4441_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_887 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_572 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5096__A _5081_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_733 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_929 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4888__A1 _4865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4888__B2 _4887_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_276 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_480 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3560__A1 _3251_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_950 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3560__B2 _3397_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_995 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3344__A _3344_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_537 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_239 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2982__B1_N _2888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4159__B _4159_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_358 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3998__B _3964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_743 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1009 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_884 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_489 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4812__A1 _4811_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_681 VGND VPWR sky130_fd_sc_hd__decap_3
X_4901_ _4900_/A _4899_/X _4900_/X _4914_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_34_843 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_342 VGND VPWR sky130_fd_sc_hd__decap_6
X_4832_ _4821_/X _4832_/B _4833_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4903__A _4914_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4025__C1 _4024_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_684 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_695 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_397 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_194 VGND VPWR sky130_fd_sc_hd__decap_12
X_4763_ _2737_/A _3875_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_712 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_403 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3519__A _3519_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4613__A2_N _4610_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_745 VGND VPWR sky130_fd_sc_hd__decap_12
X_3714_ _3713_/X _3714_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4694_ _5521_/Q _2842_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_447 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1018 VGND VPWR sky130_fd_sc_hd__fill_2
X_3645_ _5311_/Y _3644_/X _5311_/Y _3644_/X _3645_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_940 VGND VPWR sky130_fd_sc_hd__decap_12
X_3576_ _3575_/X _3600_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_804 VGND VPWR sky130_fd_sc_hd__fill_2
X_5315_ _5284_/Y _5313_/X _5350_/A _5317_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__5545__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_526 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3254__A _3305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_483 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_848 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_548 VGND VPWR sky130_fd_sc_hd__decap_12
X_5246_ _3603_/A _5245_/B _5278_/A _5246_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__4069__B _4069_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5247__B1_N _5217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_913 VGND VPWR sky130_fd_sc_hd__fill_2
X_5177_ _2696_/A _5281_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_935 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_637 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_592 VGND VPWR sky130_fd_sc_hd__decap_8
X_4128_ _4786_/X _4111_/X _4128_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_56_434 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_607 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_776 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3701__B _3689_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4059_ _4043_/C _4058_/X _4059_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_45_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_415 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_832 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_692 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_843 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_353 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_326 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4813__A _4813_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_347 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_879 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3429__A _3426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_570 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_918 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3148__B key_in[83] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_726 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_736 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_491 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_642 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_664 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_781 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_634 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3082__B1_N _3127_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4098__A2 _5540_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_986 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_66 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_166 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_881 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3845__A2 _3821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_72 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3611__B _3610_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3058__B1 _3128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_128 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_437 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_692 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2805__B1 _2814_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5418__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_312 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_367 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_520 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3230__B1 _3227_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_542 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3781__A1 _3778_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_929 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_501 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5568__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3347__A1_N _3342_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3430_ _3431_/A _3431_/B _3432_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_125_940 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3533__B2 _3532_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3361_ _3361_/A _3359_/Y _3362_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4730__B1 data_out2[26] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_910 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3074__A _3074_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_483 VGND VPWR sky130_fd_sc_hd__fill_2
X_5100_ _5473_/Q _5104_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_44_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3292_ _3293_/A key_in[23] _3292_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_345 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4089__A2 _3976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_987 VGND VPWR sky130_fd_sc_hd__decap_12
X_5031_ _5001_/X _5017_/X _5009_/X _5017_/A _5017_/B _5031_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_97_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_166 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3802__A _3795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3836__A2 _3697_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_423 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_713 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_798 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_724 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3049__B1 _3048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_990 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3915__A1_N _3058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_757 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4797__B1 data_out1[31] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_971 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_807 VGND VPWR sky130_fd_sc_hd__decap_12
X_4815_ _4815_/A _4815_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_166_317 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5210__B2 _5209_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3249__A _3248_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4746_ _4701_/A _4746_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4071__C _4784_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_4677_ _4677_/A _4677_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3628_ _3608_/X _3611_/X _3628_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_707 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5183__B key_in[32] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3524__B2 _3523_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4721__B1 data_out2[22] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_910 VGND VPWR sky130_fd_sc_hd__decap_4
X_3559_ _3396_/X _3523_/X _3526_/X _3559_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_131_932 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_280 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3415__C _3414_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_879 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5277__A1 _5253_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5229_ _5229_/A _2716_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4808__A _5448_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3827__A2 _3825_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_456 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5029__A1 _5027_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4527__B _4578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_916 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3431__B _3431_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_20 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4237__C1 _4236_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_768 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_802 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4543__A _5547_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_112 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_610 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_481 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_183 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5358__B _5357_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4262__B _4654_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_167 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5201__A1 _5199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_178 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3159__A _3182_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_189 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_339 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5201__B2 _5200_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_389 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3776__A2_N _3775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_349 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_501 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2998__A _2998_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_715 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_50 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_567 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_707 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_718 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_910 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5524__D _5524_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_87 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5268__A1 _5234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_976 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_827 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4718__A _3905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3818__A2 _3816_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1000 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_595 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_223 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4779__B1 data_out1[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_565 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3046__A3 _3041_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_971 VGND VPWR sky130_fd_sc_hd__decap_4
X_2930_ _2930_/A _2925_/Y _2930_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3995__C _3994_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4453__A _4449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_829 VGND VPWR sky130_fd_sc_hd__fill_2
X_2861_ _2861_/A key_in[75] _2861_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5390__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3069__A _3069_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4600_ _4600_/A _4600_/B _4601_/B VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2792_ _2968_/A key_in[105] _2828_/A _2792_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_12_890 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_884 VGND VPWR sky130_fd_sc_hd__fill_2
X_4531_ _4546_/A _4531_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4900__B _4899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_512 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5284__A _5515_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_394 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2701__A _3603_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_236 VGND VPWR sky130_fd_sc_hd__decap_12
X_4462_ _4469_/A _4468_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4901__B1_N _4900_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3506__A1 _5128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3516__B _3516_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_409 VGND VPWR sky130_fd_sc_hd__decap_3
X_3413_ _3340_/X _3413_/B _3413_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4393_ _4390_/X _4393_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5434__D _5434_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_610 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_280 VGND VPWR sky130_fd_sc_hd__decap_12
X_3344_ _3344_/A _3296_/X _3344_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_97_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_954 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_751 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_442 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5259__A1 _3608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5537__RESET_B _4317_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5259__B2 _5258_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_784 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4628__A _3501_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3275_ _4720_/X _3274_/X _3275_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_5014_ _4559_/A _4997_/X _5014_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_27_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_735 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3690__B1 _3681_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_532 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_554 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_587 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4363__A _4367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_598 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3869__A1_N _3866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_350 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_361 VGND VPWR sky130_fd_sc_hd__decap_4
X_4729_ _4728_/X _4725_/X data_out2[25] _4726_/X _5427_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4810__B _4810_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_523 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5194__A _3573_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3707__A _3727_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_556 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_707 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3426__B _3388_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_921 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_827 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_998 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4538__A _4537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4273__A _4271_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3433__B1 _3393_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5088__B _5086_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_963 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5519__D _5519_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_996 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3736__A1 _3726_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_670 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_168 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_60 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2704__B1_N _2686_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_692 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3617__A _3600_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_707 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_504 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5313__A1_N _5286_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3336__B key_in[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_418 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4161__A1 _4128_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_602 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4448__A _4469_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_326 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2894__C _2821_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_646 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3352__A _3284_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_123 VGND VPWR sky130_fd_sc_hd__fill_1
X_3060_ _3060_/A _3060_/B _3060_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_979 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4167__B _4090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3071__B _3071_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_521 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_863 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_351 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5279__A _5277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_587 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4183__A _4092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_738 VGND VPWR sky130_fd_sc_hd__fill_2
X_3962_ _3959_/X _3961_/Y _3962_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_44_790 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4614__C _4614_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_952 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3975__A1 data_in1[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_615 VGND VPWR sky130_fd_sc_hd__fill_2
X_2913_ _2913_/A _2912_/X _2913_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_148_103 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4599__A1_N _4600_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5429__D _4732_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3893_ _3886_/X _3892_/X _3893_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_149_659 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4911__A _4911_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2844_ _2855_/A _2844_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_148_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_629 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4924__B1 _5554_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_670 VGND VPWR sky130_fd_sc_hd__fill_1
X_5563_ _4562_/X _5563_/Q _4287_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2775_ _2735_/X _2774_/B _2784_/A _2778_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3606__A2_N _3605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_320 VGND VPWR sky130_fd_sc_hd__fill_1
X_4514_ _4515_/A _4514_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_545 VGND VPWR sky130_fd_sc_hd__decap_4
X_5494_ _5494_/D _5494_/Q _4370_/X _5430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_813 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_578 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_206 VGND VPWR sky130_fd_sc_hd__decap_8
X_4445_ _4443_/A _4445_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_172_695 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_4376_ _4397_/A _4381_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_985 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5371__RESET_B _4515_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_913 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4358__A _4354_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3327_ _3155_/Y _3324_/B _3326_/Y _3331_/A VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_112_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_935 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3262__A _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_3258_ _3258_/A _3258_/B _3258_/C _3258_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_85_156 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4077__B _4076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_49 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_39 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_584 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_329 VGND VPWR sky130_fd_sc_hd__fill_2
X_3189_ _3145_/X key_in[52] _3189_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_9 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_223 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_757 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_768 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5189__A _4798_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4093__A _4074_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_952 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_37 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_935 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_782 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4821__A _4821_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_495 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3718__A1 data_in1[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4540__B _4541_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3437__A _3419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_556 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_30 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5459__RESET_B _4411_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_812 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2941__A2 _5497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_846 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_323 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_183 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4143__A1 data_in1[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_345 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5340__B1 _5338_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_602 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3449__B1_N _3416_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_473 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4268__A _4267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3172__A _5222_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3900__A _3835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_576 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_384 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_259 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_985 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_434 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4731__A _5538_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_467 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3709__B2 _3708_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4906__B1 _4905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_810 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_843 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3066__B _3066_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_813 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3592__A2_N _3591_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4230_ _4794_/X _4212_/X _4230_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_141_367 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4685__A2 _4674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5281__B _5281_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4161_ _4128_/X _4160_/X _4138_/X _4198_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__4178__A _4791_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_3112_ _3038_/A _3112_/B _3037_/Y _3112_/X VGND VPWR sky130_fd_sc_hd__or3_4
X_4092_ _3569_/A _4092_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_3043_ _2859_/A _3043_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3645__B1 _5311_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_830 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_513 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_693 VGND VPWR sky130_fd_sc_hd__decap_12
X_4994_ _4896_/X _4991_/Y _4992_/X _4993_/Y _4806_/X _5464_/D VGND VPWR sky130_fd_sc_hd__a32oi_4
XANTENNA__3948__A1 data_in1[17] VGND VPWR sky130_fd_sc_hd__diode_2
X_3945_ _3945_/A _3945_/B _3945_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4070__B1 _4043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_911 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_281 VGND VPWR sky130_fd_sc_hd__fill_2
X_3876_ _3826_/Y _3875_/X _3851_/X _3876_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_149_478 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_618 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_489 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_810 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_949 VGND VPWR sky130_fd_sc_hd__fill_2
X_2827_ _2898_/A _2859_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_136_128 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3257__A _3187_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5175__C _3573_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5546_ _4542_/X _4542_/A _4307_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2758_ _4637_/A _2754_/X _2755_/X _2756_/X _2757_/X _2759_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_117_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5552__RESET_B _4300_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_802 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_824 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_5477_ _5477_/D _5477_/Q _4389_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2689_ _2687_/X _2688_/X _2687_/X _2688_/X _2689_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_4428_ _4426_/X _4428_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_120_507 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3704__B _3703_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_15 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4088__A _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2687__A1 _4859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1006 VGND VPWR sky130_fd_sc_hd__fill_1
X_4359_ _4354_/X _4359_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_690 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_87 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4535__B _4542_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_58 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_716 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_587 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_896 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_822 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_524 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_749 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_535 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_248 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4551__A _5554_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_242 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_776 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5451__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_916 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_904 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_977 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5366__B key_in[38] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_414 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_297 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_448 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3167__A2 _3166_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_95 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_375 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2914__A2 _2912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_621 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4116__A1 _4784_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_99 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5313__B1 _5286_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_507 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5532__D _5532_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_104 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3623__A1_N _5272_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4726__A _4701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_446 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3630__A _3630_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_852 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_479 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_844 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_888 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4052__B1 _4051_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4461__A _4461_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3730_ _3730_/A _3730_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_60_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_765 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_927 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5276__B _5276_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_629 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_286 VGND VPWR sky130_fd_sc_hd__decap_12
X_3661_ _3660_/X _3661_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4180__B _4196_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5191__A1_N _5182_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_448 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3077__A _3077_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5400_ _4796_/X data_out1[30] _4481_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_146_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VPWR sky130_fd_sc_hd__decap_8
X_3592_ _5213_/X _3591_/X _5213_/X _3591_/X _3592_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_115_802 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_684 VGND VPWR sky130_fd_sc_hd__fill_1
X_5331_ _5331_/A _5332_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_47_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_846 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_492 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_480 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5292__A _5262_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3805__A _3804_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5304__B1 _2828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_345 VGND VPWR sky130_fd_sc_hd__decap_4
X_5262_ _3626_/A _5262_/B _5262_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_687 VGND VPWR sky130_fd_sc_hd__decap_12
X_4213_ _4794_/X _4212_/X _4213_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_849 VGND VPWR sky130_fd_sc_hd__decap_4
X_5193_ _5198_/B _5226_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5442__D _4599_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_432 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3866__B1 _2980_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_808 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3330__A2 _3328_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_977 VGND VPWR sky130_fd_sc_hd__decap_4
X_4144_ _4126_/X _4090_/X _3231_/A _4144_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_56_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_796 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_4075_ _4073_/X _4074_/X _4075_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__4636__A _4636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3540__A _3540_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5083__A2 _5079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_148 VGND VPWR sky130_fd_sc_hd__decap_12
X_3026_ _3026_/A _2884_/B _5527_/Q _3026_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_71_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_800 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3094__B2 _3093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_980 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_682 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4228__A2_N _4227_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_129 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2841__B2 _2840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5474__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_877 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4977_ _4997_/C _4976_/X _4997_/C _4976_/X _4978_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4371__A _4375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3928_ data_in1[16] _3837_/X _3902_/X _3927_/Y _3928_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_149_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_16 VGND VPWR sky130_fd_sc_hd__decap_4
X_3859_ _3769_/Y _5530_/Q _2842_/A _3858_/Y _3859_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_137_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_768 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3149__A2 key_in[115] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_960 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_418 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_982 VGND VPWR sky130_fd_sc_hd__fill_2
X_5529_ _3142_/X _5529_/Q _4328_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_3_428 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3715__A _3712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_367 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3434__B _3364_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_197 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_329 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_958 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4546__A _4546_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3450__A _3450_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_852 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5074__A2 _5072_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_502 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_844 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_630 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_855 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_96 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__B1 _3230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_899 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_538 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4281__A _4276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_916 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5474__RESET_B _4393_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5096__B _5096_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_701 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_949 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_774 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5527__D _5527_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5403__RESET_B _4478_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_778 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4888__A2 _4877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_183 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3625__A _3618_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_440 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3560__A2 _5510_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_985 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_462 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3344__B _3296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_483 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4159__C _4120_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_605 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_733 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4456__A _4461_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3998__C _3952_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3360__A _3361_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_852 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5497__CLK _5429_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_243 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4812__A2 _4810_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_287 VGND VPWR sky130_fd_sc_hd__decap_12
X_4900_ _4900_/A _4899_/X _4900_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2823__A1 _2822_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4831_ _4830_/A _4830_/B _4830_/X _4833_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__4025__B1 _3997_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4903__B _4902_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_162 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5287__A _5287_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4191__A _4189_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4762_ _2714_/A _4757_/X data_out1[12] _4758_/X _5382_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_159_562 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1005 VGND VPWR sky130_fd_sc_hd__fill_2
X_3713_ _4750_/X _3690_/X _3693_/X _3713_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3519__B _2885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_415 VGND VPWR sky130_fd_sc_hd__decap_12
X_4693_ _2847_/A _4687_/X data_out2[9] _4688_/X _5411_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__5437__D _5437_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_3644_ _3641_/A _3640_/X _3666_/B _3644_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_128_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_3575_ _5190_/Y _3574_/X _5190_/Y _3574_/X _3575_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_952 VGND VPWR sky130_fd_sc_hd__decap_6
X_5314_ _5284_/Y _5313_/X _5350_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_451 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_996 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2771__A1_N _2762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5245_ _3603_/A _5245_/B _5278_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_197 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4069__C _4069_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_903 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_605 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_5176_ _5355_/A _2696_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_69_785 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_104 VGND VPWR sky130_fd_sc_hd__fill_1
X_4127_ _4126_/X _4090_/X _4788_/X _4127_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_29_649 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4366__A _4367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3270__A _3227_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_468 VGND VPWR sky130_fd_sc_hd__decap_12
X_4058_ _4046_/Y _4057_/X _4046_/Y _4057_/X _4058_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_619 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_3009_ _3050_/B _3008_/Y _3050_/B _3008_/Y _3892_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_855 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_305 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_315 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_316 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_140 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4813__B _4812_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5197__A _5197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3429__B _3429_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_554 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_565 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_971 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_470 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_790 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_930 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_748 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3445__A _3501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_943 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_936 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_50 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4276__A _4304_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_40 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3180__A _3180_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_84 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3058__B2 _3057_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2805__B2 _2804_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_641 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_866 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_961 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_983 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_893 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_724 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3230__B2 _3229_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_520 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_908 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_554 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3781__A2 _3777_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_418 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3518__C1 _3517_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_952 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4245__A1_N _4239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4730__A1 _5537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3360_ _3361_/A _3359_/Y _3362_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_125_985 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_825 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4730__B2 _4726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_922 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3074__B _3071_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_313 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_270 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_495 VGND VPWR sky130_fd_sc_hd__fill_2
X_3291_ _3291_/A key_in[55] _3291_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_292 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_808 VGND VPWR sky130_fd_sc_hd__decap_12
X_5030_ _5034_/A _5030_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_25_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_999 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3297__A1 _5470_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_925 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3802__B _3801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4186__A _4170_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_435 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3090__A _3090_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3049__A1 _5463_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_660 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4797__A1 _5510_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4914__A _4886_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4797__B2 _4677_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_19 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5396__RESET_B _4486_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_983 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_825 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_471 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_819 VGND VPWR sky130_fd_sc_hd__decap_12
X_4814_ _4813_/A _4812_/X _4814_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_33_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_493 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3249__B _3249_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_381 VGND VPWR sky130_fd_sc_hd__decap_4
X_4745_ _4699_/A _4745_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_21_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5512__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_908 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_245 VGND VPWR sky130_fd_sc_hd__decap_4
X_4676_ _4700_/A _4677_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3454__A1_N _3438_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_598 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_3627_ _3626_/A _3625_/X _3626_/X _3630_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_89_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4721__A1 _4720_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3558_ _3522_/X _3536_/X _4661_/X _3562_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4721__B2 _4713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_292 VGND VPWR sky130_fd_sc_hd__decap_4
X_3489_ _3489_/A _3541_/C _3491_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5277__A2 _5276_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_977 VGND VPWR sky130_fd_sc_hd__decap_4
X_5228_ _5481_/Q _3608_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_57_700 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_571 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_722 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4096__A _4095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_733 VGND VPWR sky130_fd_sc_hd__fill_2
X_5159_ _5159_/A _5159_/B _5160_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__5029__A2 _5027_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4527__C _4525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_928 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4237__B1 _4221_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_276 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_585 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4824__A _4822_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_961 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_268 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3996__C1 _3995_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_279 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4543__B _4542_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_58 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_313 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_493 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_146 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5201__A2 _5361_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_317 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3159__B _3159_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_863 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2998__B _2998_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2971__B1 _2828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3175__A _3175_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_545 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_952 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_421 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3903__A _3884_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_99 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5268__A2 key_in[99] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5540__D _3518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_541 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_788 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4228__B1 _4222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4779__A1 _4778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_758 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4734__A _5540_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4779__B2 _4770_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_909 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_235 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_674 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3451__A1 _3450_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_983 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_791 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5535__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_493 VGND VPWR sky130_fd_sc_hd__decap_12
X_2860_ _2861_/A key_in[11] _2860_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3069__B _3068_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5246__B1_N _5278_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_880 VGND VPWR sky130_fd_sc_hd__decap_4
X_2791_ _2898_/A _2968_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_157_852 VGND VPWR sky130_fd_sc_hd__fill_2
X_4530_ _4529_/X _4546_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_172_800 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_42 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_738 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_4461_ _4461_/A _4461_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_7_86 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3085__A _3085_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_248 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_3412_ _5472_/Q _3379_/B _3412_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3506__A2 _3474_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4392_ _4390_/X _4392_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_590 VGND VPWR sky130_fd_sc_hd__decap_12
X_3343_ _5470_/Q _3295_/X _3343_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4909__A _4873_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_966 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3813__A _3569_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5259__A2 _2717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_666 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_454 VGND VPWR sky130_fd_sc_hd__decap_4
X_3274_ _3250_/Y _3273_/X _3250_/Y _3273_/X _3274_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_999 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_796 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_5013_ _5013_/A _5017_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5450__D _4835_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_541 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_777 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_703 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5577__RESET_B _4270_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_928 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_725 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3690__B2 _3689_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5506__RESET_B _4355_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_758 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4644__A _4522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3442__A1 _3441_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4137__A1_N _4130_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_791 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_17 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_655 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_627 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_104 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_137 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_699 VGND VPWR sky130_fd_sc_hd__decap_3
X_2989_ _2989_/A _2989_/B _2989_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4728_ _5536_/Q _4728_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_162_310 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3707__B _3687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5194__B _5226_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_4659_ _4576_/X _4666_/D _4658_/X _4659_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_162_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_343 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3426__C _3359_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_899 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_933 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_537 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4819__A _4819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_655 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3723__A _2735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5408__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_98 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_699 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_349 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_917 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3130__B1 _3125_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_596 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5558__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_544 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4554__A _4554_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_769 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_728 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3433__A1 data_in2[26] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_830 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_147 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3736__A2 _3733_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2802__A _2802_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_118 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_810 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_72 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3617__B _3616_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_832 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_843 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5535__D _3363_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_866 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_760 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_887 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4697__B1 data_out2[11] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4161__A2 _4160_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_752 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3633__A _3615_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_817 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_925 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3352__B _3352_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5110__A1 _5090_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_338 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4167__C _4791_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_552 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3121__B1 _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3071__C _3071_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_308 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3672__A1 _3671_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_736 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_831 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4464__A _4468_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_235 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5279__B _5280_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_363 VGND VPWR sky130_fd_sc_hd__decap_12
X_3961_ _3908_/Y _3935_/X _3960_/X _3961_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__4183__B _4183_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_599 VGND VPWR sky130_fd_sc_hd__fill_2
X_2912_ _2910_/Y _2911_/X _2912_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3975__A2 _3837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_964 VGND VPWR sky130_fd_sc_hd__decap_12
X_3892_ _3892_/A _3891_/X _3892_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_31_463 VGND VPWR sky130_fd_sc_hd__decap_12
X_2843_ _2842_/X _2855_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4911__B _4910_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5295__A _5294_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3808__A _3791_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2712__A _2770_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5562_ _4561_/X _5562_/Q _4288_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_163_107 VGND VPWR sky130_fd_sc_hd__decap_3
X_2774_ _2735_/X _2774_/B _2784_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4924__B2 _4923_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_822 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2935__B1 _2828_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4513_ _4515_/A _4513_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_156_192 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5445__D _4612_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5493_ _5493_/D _2797_/A _4371_/X _5430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_172_652 VGND VPWR sky130_fd_sc_hd__decap_12
X_4444_ _4443_/A _4444_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_825 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3130__A2_N _3129_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4639__A _4638_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4375_ _4375_/A _4375_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3543__A _3543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_903 VGND VPWR sky130_fd_sc_hd__decap_4
X_3326_ _3325_/X _3326_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_997 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_785 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_593 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3262__B key_in[22] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_647 VGND VPWR sky130_fd_sc_hd__decap_12
X_3257_ _3187_/A _3257_/B _3186_/Y _3258_/C VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_74_809 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_168 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_883 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_clock clkbuf_3_7_0_clock/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_54_511 VGND VPWR sky130_fd_sc_hd__decap_8
X_3188_ _3187_/A _3186_/Y _3187_/X _3188_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_82_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_842 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4374__A _4375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5189__B _5189_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_16 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4093__B _4082_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4612__B1 _4611_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_238 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_430 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_947 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4821__B _4821_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_457 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3179__B1 _3902_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4915__A1 _4900_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3718__A2 _3697_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_669 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_513 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3437__B _3419_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_140 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_814 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_195 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4143__A2 _4125_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5340__A1 _4636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4549__A _5552_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5340__B2 _5339_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_357 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_752 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5499__RESET_B _4364_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3351__B1 _3316_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5428__RESET_B _4449_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5380__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_628 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_56 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_725 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_127 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4851__B1 _5548_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3900__B _3898_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4284__A _4289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_588 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_599 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_536 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_794 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4915__B1_N _4914_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3628__A _3608_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4906__A1 _4896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_660 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4906__B2 _4806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_682 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2917__B1 _2888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_833 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_855 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_343 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3590__B1 _4679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_376 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4459__A _4461_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_346 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3238__A1_N _3230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3342__B1 _3341_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5281__C _5281_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4160_ _4788_/X _4137_/X _4160_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4178__B _4177_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_3111_ _3110_/A _3110_/B _3160_/A _3116_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_67_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_744 VGND VPWR sky130_fd_sc_hd__fill_2
X_4091_ _4026_/A _4090_/X _4786_/X _4091_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5095__B1 _5109_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3042_ _2861_/A key_in[80] _3042_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_788 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3645__B2 _3644_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_691 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4194__A _3466_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2707__A _2707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2853__C1 _2852_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_672 VGND VPWR sky130_fd_sc_hd__fill_2
X_4993_ _4985_/X _4993_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_23_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_536 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4922__A _5553_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1003 VGND VPWR sky130_fd_sc_hd__decap_12
X_3944_ _2889_/Y _3941_/X _3943_/X _3945_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3948__A2 _3837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4070__A1 data_in1[22] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_569 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_794 VGND VPWR sky130_fd_sc_hd__fill_1
X_3875_ _3875_/A _3850_/X _3875_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_104_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_608 VGND VPWR sky130_fd_sc_hd__fill_2
X_2826_ _2861_/A key_in[74] _2826_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_158_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_833 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3257__B _3257_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5545_ _4541_/X _4541_/A _4308_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_641 VGND VPWR sky130_fd_sc_hd__fill_1
X_2757_ _5300_/A key_in[104] _2828_/A _2757_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_118_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_5476_ _5476_/D _5143_/A _4391_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_696 VGND VPWR sky130_fd_sc_hd__fill_1
X_2688_ _5335_/X _2769_/A _5343_/X _2688_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_133_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_633 VGND VPWR sky130_fd_sc_hd__decap_8
X_4427_ _4426_/X _4427_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4369__A _4397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3273__A _3273_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3333__B1 _3332_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4358_ _4354_/X _4358_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_783 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3084__A2_N _3083_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2687__A2 _2686_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4088__B _4088_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_794 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5521__RESET_B _4337_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_733 VGND VPWR sky130_fd_sc_hd__decap_6
X_3309_ _3287_/C _3309_/B _3309_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_171_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_444 VGND VPWR sky130_fd_sc_hd__decap_12
X_4289_ _4289_/A _4289_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_232 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5086__B1 _5084_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_864 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_599 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5312__A1_N _5297_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_32 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4832__A _4821_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_14 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_65 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_733 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_772 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_36 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4551__B _4547_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_934 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_989 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_426 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_490 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_961 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_343 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_983 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_888 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_825 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_471 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4116__A2 _4083_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4279__A _4276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5313__B2 _5322_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_654 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3183__A _3116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_219 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_699 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_187 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_967 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3911__A _3861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3627__A1 _3626_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3605__A2_N _3604_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3630__B _3628_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_190 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_352 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_525 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4052__A1 _3932_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_366 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_591 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3358__A _3210_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3162__A1_N _3154_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_939 VGND VPWR sky130_fd_sc_hd__decap_12
X_3660_ _5516_/Q _3659_/X _3660_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_158_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_427 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3077__B key_in[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_3591_ _3573_/X _3590_/X _3573_/X _3590_/X _3591_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_419 VGND VPWR sky130_fd_sc_hd__decap_8
X_5330_ _5330_/A _5331_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3563__B1 _3557_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_696 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3805__B _3803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_121 VGND VPWR sky130_fd_sc_hd__fill_1
X_5261_ _5261_/A _5262_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5304__A1 _5300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_132 VGND VPWR sky130_fd_sc_hd__decap_12
X_4212_ _4212_/A _4211_/X _4212_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_69_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_176 VGND VPWR sky130_fd_sc_hd__fill_2
X_5192_ _5178_/Y _5198_/B _5192_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_123_891 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_945 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3866__B2 _3865_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4143_ data_in1[25] _4125_/X _4127_/X _4142_/Y _4143_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4917__A _4917_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_904 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3821__A _3799_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_403 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_786 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_105 VGND VPWR sky130_fd_sc_hd__decap_8
X_4074_ _4045_/X _4057_/X _4074_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_499 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_585 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_959 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3540__B _3540_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3025_ data_in2[15] _2956_/X _2996_/X _3024_/Y _3025_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_93_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_322 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_193 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4652__A _4819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5240__B1 _5211_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4976_ _4555_/A _4965_/X _4975_/X _4976_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3927_ _3835_/A _3925_/Y _3926_/X _3927_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_3858_ _5530_/Q _3858_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_20_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_2809_ _2784_/Y _2846_/B _2809_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_118_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_246 VGND VPWR sky130_fd_sc_hd__decap_6
X_3789_ data_in1[10] _3697_/X _3765_/X _3788_/Y _3789_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3554__B1 _3552_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2900__A _2790_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5528_ _3101_/X _5528_/Q _4329_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_146_994 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_173 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_493 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_324 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_121 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3715__B _3714_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_964 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4099__A _3980_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5459_ _4941_/X _4642_/A _4411_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_121_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3306__B1 _3304_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3434__C _4731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_742 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4827__A _4827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_775 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_477 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_820 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3609__A1 _3608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_596 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3450__B _3449_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_352 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_812 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_897 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_672 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_311 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4562__A _5563_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3591__A2_N _3590_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_664 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__B2 _4033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5231__B1 _5230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3178__A _3178_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_747 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_724 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_786 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_746 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_950 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4888__A3 _4866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_600 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_267 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2810__A _2852_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_493 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_633 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5443__RESET_B _4430_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_930 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3625__B _3624_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_195 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_290 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5543__D _5543_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_132 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_963 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_496 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_764 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4737__A _4701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_861 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3641__A _3641_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_797 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_285 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3998__D _3987_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_436 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_831 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_296 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3360__B _3359_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_469 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_650 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_299 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_631 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2823__A2 _2821_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_653 VGND VPWR sky130_fd_sc_hd__decap_12
X_4830_ _4830_/A _4830_/B _4830_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4472__A _4475_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_355 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4025__A1 data_in1[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_517 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_174 VGND VPWR sky130_fd_sc_hd__decap_4
X_4761_ _3804_/A _4757_/X data_out1[11] _4758_/X _4761_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_21_539 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4191__B _4190_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3088__A _2889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3784__B1 _3759_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3712_ _2717_/A _3710_/X _3741_/A _3712_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_147_725 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3519__C _5541_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4692_ _5520_/Q _2847_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_3643_ _3642_/X _3666_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_128_983 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3536__B1 _3527_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_780 VGND VPWR sky130_fd_sc_hd__fill_2
X_3574_ _5178_/Y _3572_/Y _3573_/X _3574_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_115_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_622 VGND VPWR sky130_fd_sc_hd__fill_2
X_5313_ _5286_/Y _5322_/A _5286_/Y _5322_/A _5313_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5453__D _4869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_964 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_441 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5289__B1 _3577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_5244_ _5227_/Y _5243_/X _5227_/Y _5243_/X _5245_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4116__B1_N _4115_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5175_ _5197_/A _5252_/B _3573_/A _5175_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3551__A _3529_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_712 VGND VPWR sky130_fd_sc_hd__decap_12
X_4126_ _4537_/X _4126_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5441__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_425 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_948 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_894 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_222 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3270__B _3269_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4057_ _3273_/B _4056_/X _3273_/B _4056_/X _4057_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3008_ _2974_/Y _2978_/X _2973_/Y _3008_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_71_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_642 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_867 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4382__A _4381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_317 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_45 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_339 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_377 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5197__B _5252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_38 VGND VPWR sky130_fd_sc_hd__fill_2
X_4959_ _4954_/Y _4958_/B _4958_/X _4961_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_138_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_500 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_599 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_482 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3445__B key_in[91] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_603 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_955 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_658 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4557__A _4997_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_296 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3180__B _3180_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_907 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_970 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4292__A _4296_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_303 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_94 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_174 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_848 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3215__C1 _3214_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5538__D _5538_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_347 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_9 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_500 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_511 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_717 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3636__A _5520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3518__B1 _3493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_964 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4730__A2 _4725_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_761 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4227__A2_N _4226_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5464__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_782 VGND VPWR sky130_fd_sc_hd__decap_8
X_3290_ _4582_/X _3318_/A _3290_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_151_282 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_292 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4467__A _4468_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_509 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3297__A2 _3295_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_937 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4186__B _4176_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_959 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_691 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3090__B _3038_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_918 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3049__A2 _3047_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_428 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3498__A2_N _3497_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4914__B _4914_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4797__A2 _4674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5298__A _5234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_995 VGND VPWR sky130_fd_sc_hd__decap_12
X_4813_ _4813_/A _4812_/X _4823_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3421__A2_N _3420_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5448__D _4816_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_347 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3757__B1 _3720_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4930__A _4815_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3249__C _3176_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_371 VGND VPWR sky130_fd_sc_hd__fill_1
X_4744_ _5260_/A _4736_/X data_out1[3] _4737_/X _5373_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_119_224 VGND VPWR sky130_fd_sc_hd__decap_3
X_4675_ _4672_/X _4700_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3509__B1 _3498_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3626_ _3626_/A _3625_/X _3626_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_3557_ _3548_/Y _3556_/Y _3548_/Y _3556_/Y _3557_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4721__A2 _4712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_452 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_975 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2692__A2_N _2691_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_945 VGND VPWR sky130_fd_sc_hd__decap_4
X_3488_ _3488_/A _3488_/B _3488_/C _3487_/Y _3541_/C VGND VPWR sky130_fd_sc_hd__nor4_4
X_5227_ _5256_/A _5227_/B _5227_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_103_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_455 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4377__A _4381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_550 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_168 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_712 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_892 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_5158_ _5159_/A _5159_/B _5160_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_56_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_391 VGND VPWR sky130_fd_sc_hd__decap_6
X_4109_ _3347_/X _4108_/Y _3347_/X _4108_/Y _4109_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_767 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4527__D _4629_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_5089_ _4870_/X _5087_/Y _5096_/B _5076_/A _4930_/X _5089_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4237__A1 data_in1[30] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_203 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_480 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4824__B _4825_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_631 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3996__B1 _3978_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_973 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5001__A _5001_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_809 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_136 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_325 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_147 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_319 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4840__A _4840_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_831 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_881 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_544 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_380 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_886 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2998__C _2998_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3456__A _4731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2971__A1 _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_739 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5487__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_780 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_964 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_956 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3903__B _3893_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4287__A _4289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_509 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3191__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_51 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_84 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_704 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_266 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4228__B2 _4227_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_428 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4779__A2 _4769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3987__B1 _3154_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3451__A2 _3449_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_133 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4151__A2_N _4150_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4750__A _5200_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ _2790_/A key_in[73] _2790_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_864 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_380 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3366__A _3366_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2962__A1 _2961_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4460_ _4461_/A _4460_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_227 VGND VPWR sky130_fd_sc_hd__decap_6
X_3411_ _5473_/Q _3410_/X _5473_/Q _3410_/X _3416_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_290 VGND VPWR sky130_fd_sc_hd__fill_2
X_4391_ _4390_/X _4391_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_125_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_3342_ _5076_/A _3340_/B _3341_/Y _3342_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_97_111 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_731 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4909__B _4908_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4197__A _4158_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3273_ _3273_/A _3273_/B _3273_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_85_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_689 VGND VPWR sky130_fd_sc_hd__decap_12
X_5012_ _4996_/A _4995_/X _4942_/X _5011_/Y _5012_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_66_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_907 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_553 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_873 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4925__A _4925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_288 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4644__B _4576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_940 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_962 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_601 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3442__A2 _3441_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_921 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5546__RESET_B _4307_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_100 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1004 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3990__A2_N _3989_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_116 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4660__A _5256_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_818 VGND VPWR sky130_fd_sc_hd__fill_2
X_2988_ _2925_/A _2988_/B _2924_/Y _2988_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_21_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_864 VGND VPWR sky130_fd_sc_hd__decap_12
X_4727_ _3316_/C _4725_/X data_out2[24] _4726_/X _5426_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_148_886 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_10_0_clock clkbuf_3_5_0_clock/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3276__A _3275_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_823 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_300 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_845 VGND VPWR sky130_fd_sc_hd__fill_2
X_4658_ _4525_/X _4586_/B _4519_/X _4253_/D _4658_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_135_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_867 VGND VPWR sky130_fd_sc_hd__decap_8
X_3609_ _3608_/A _3607_/X _3608_/X _3609_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_163_889 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_506 VGND VPWR sky130_fd_sc_hd__decap_12
X_4589_ _4589_/A _4588_/Y _4590_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_103_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_783 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_945 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4819__B _4818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_293 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3723__B _3722_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_764 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_818 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_851 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3130__B2 _3129_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_361 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_586 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_737 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4554__B _4547_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_984 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_461 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_601 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3433__A2 _3391_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_617 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4570__A _5129_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_352 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2802__B _2801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3186__A _3159_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_855 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_878 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4697__A1 _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_208 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_772 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_219 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4697__B2 _4688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_398 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_72 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3633__B _3570_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5551__D _4548_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_571 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5110__A2 _5093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_199 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_840 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3121__A1 _3043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_158 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5502__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4745__A _4699_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_501 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_884 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3672__A2 _3670_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3453__A1_N _3442_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_748 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_394 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_843 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_876 VGND VPWR sky130_fd_sc_hd__decap_8
X_3960_ _3073_/C _3935_/B _3960_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_898 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4183__C _4183_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2911_ _2838_/A _2865_/X _2834_/X _2770_/Y _2911_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_3891_ _3890_/X _3891_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_43_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_976 VGND VPWR sky130_fd_sc_hd__fill_1
X_2842_ _2842_/A _2842_/B _2842_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4480__A _4477_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3188__A1 _3187_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_650 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3808__B _3806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2712__B _2711_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2773_ _2736_/Y _2772_/X _2736_/Y _2772_/X _2774_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5561_ _4559_/X _4559_/A _4289_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_129_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3096__A _3073_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2935__A1 _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_160 VGND VPWR sky130_fd_sc_hd__fill_1
X_4512_ _4515_/A _4512_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_845 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_682 VGND VPWR sky130_fd_sc_hd__decap_12
X_5492_ _5492_/D _2737_/A _4372_/X _5430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_867 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4137__B1 _4130_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_664 VGND VPWR sky130_fd_sc_hd__decap_12
X_4443_ _4443_/A _4443_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3824__A _3823_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_528 VGND VPWR sky130_fd_sc_hd__fill_2
X_4374_ _4375_/A _4374_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_943 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3543__B _3543_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3325_ _3324_/X _3325_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5461__D _5461_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_241 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_615 VGND VPWR sky130_fd_sc_hd__fill_2
X_3256_ _3236_/A _3233_/X _3258_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_39_531 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_542 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4655__A _4809_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_715 VGND VPWR sky130_fd_sc_hd__fill_2
X_3187_ _3187_/A _3186_/Y _3187_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_895 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_331 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1009 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_876 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_206 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4612__A1 _4646_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_39 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5380__RESET_B _4505_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4058__A2_N _4057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_397 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_420 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_116 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4390__A _4397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2903__A _4642_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3179__A1 _3032_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_469 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3179__B2 _3178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4915__A2 _4913_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3437__C _3319_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_867 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3734__A _3726_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_36 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_420 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_720 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5340__A2 _5336_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4549__B _4541_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5525__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3351__B2 _3365_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_306 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5371__D _5371_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_873 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4565__A _5566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_512 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_981 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4851__B2 _4850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_737 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_523 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5468__RESET_B _4400_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3900__C _3899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2862__B1 _2828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_959 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2813__A _2772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_250 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_94 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_72 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3628__B _3611_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5546__D _4542_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4906__A2 _4903_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_479 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_300 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2917__B2 _2916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_630 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3590__A1 _3588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_355 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3590__B2 _5517_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_685 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_173 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_591 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3342__A1 _5076_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4136__A1_N _3382_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_881 VGND VPWR sky130_fd_sc_hd__decap_4
X_3110_ _3110_/A _3110_/B _3160_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_4090_ _4664_/X _4090_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_1_891 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5095__A1 _5090_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_467 VGND VPWR sky130_fd_sc_hd__fill_2
X_3041_ _2861_/A key_in[16] _3041_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4475__A _4475_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_821 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2853__B1 _2812_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4194__B _4193_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2707__B key_in[71] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_342 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_651 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_217 VGND VPWR sky130_fd_sc_hd__fill_2
X_4992_ _4992_/A _4990_/X _4992_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_17_792 VGND VPWR sky130_fd_sc_hd__fill_1
X_3943_ _3113_/A _3942_/Y _3943_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4922__B _4908_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4070__A2 _3976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1015 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3819__A _3819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2723__A _2723_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_935 VGND VPWR sky130_fd_sc_hd__decap_8
X_3874_ _3827_/X _3852_/X _3832_/Y _3874_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_165_907 VGND VPWR sky130_fd_sc_hd__fill_2
X_2825_ _2934_/A key_in[10] _2825_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_136_108 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5456__D _4906_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3257__C _3186_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5544_ _4540_/X _4837_/B _4309_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_129_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_845 VGND VPWR sky130_fd_sc_hd__decap_8
X_2756_ _5301_/A key_in[72] _2756_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_129_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_653 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5548__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2687_ _4859_/A _2686_/B _2686_/Y _2687_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_5475_ _5142_/X _5128_/A _4392_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_144_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_623 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_848 VGND VPWR sky130_fd_sc_hd__decap_6
X_4426_ _4419_/A _4426_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3333__A1 _3331_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3273__B _3273_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_4357_ _4354_/X _4357_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_924 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4088__C _4087_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_412 VGND VPWR sky130_fd_sc_hd__decap_12
X_3308_ _3290_/Y _3318_/B _3290_/Y _3318_/B _3309_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_594 VGND VPWR sky130_fd_sc_hd__fill_1
X_4288_ _4289_/A _4288_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_101_745 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5086__A1 _5059_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_456 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5086__B2 _5085_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_244 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_350 VGND VPWR sky130_fd_sc_hd__decap_12
X_3239_ _4661_/X _3201_/X _3177_/Y _3239_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4385__A _4387_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_255 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3097__B1 _3096_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_810 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5561__RESET_B _4289_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_320 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_876 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_887 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_695 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4832__B _4832_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_712 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3729__A _3728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_26 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_946 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_31 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_929 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_928 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_631 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_438 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_355 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3464__A _3464_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3183__B _3183_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_147 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3911__B _3891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_478 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2808__A _2784_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_489 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4295__A _4296_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_501 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_821 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3627__A2 _3625_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_832 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_556 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_567 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4052__A2 _4048_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_210 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_907 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_244 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3358__B _3357_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_294 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_406 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_254 VGND VPWR sky130_fd_sc_hd__decap_12
X_3590_ _3588_/Y _3589_/Y _4679_/X _5517_/Q _3590_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_127_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_972 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3563__B2 _3562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3374__A _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_174 VGND VPWR sky130_fd_sc_hd__decap_12
X_5260_ _5260_/A _3626_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5304__A2 key_in[100] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4211_ _3508_/X _4210_/X _3508_/X _4210_/X _4211_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5191_ _5182_/X _5190_/Y _5182_/X _5190_/Y _5198_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_924 VGND VPWR sky130_fd_sc_hd__fill_2
X_4142_ _4092_/X _4142_/B _4142_/C _4142_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_110_520 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4917__B _4915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_916 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3821__B _3819_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4073_ _3939_/X _4073_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_415 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2718__A _2718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3079__B1 _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3024_ _2927_/A _3022_/Y _3023_/X _3024_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_83_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_191 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_971 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_364 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4933__A _4921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_161 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_509 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_334 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4643__A1_N _4616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_356 VGND VPWR sky130_fd_sc_hd__decap_8
X_4975_ _4921_/X _4975_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5240__A1 _4811_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_200 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_367 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_222 VGND VPWR sky130_fd_sc_hd__fill_2
X_3926_ _3925_/A _3924_/Y _3926_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_149_233 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_581 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2983__A2_N _2982_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_592 VGND VPWR sky130_fd_sc_hd__decap_12
X_3857_ _3839_/A _3812_/B _3870_/A _3857_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5370__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_428 VGND VPWR sky130_fd_sc_hd__decap_6
X_2808_ _2784_/Y _2846_/B _2808_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3003__B1 _2828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_940 VGND VPWR sky130_fd_sc_hd__decap_6
X_3788_ _3788_/A _3786_/Y _3787_/X _3788_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_118_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3554__A1 _4640_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_804 VGND VPWR sky130_fd_sc_hd__decap_12
X_5527_ _5527_/D _5527_/Q _4330_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4751__B1 data_out1[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3554__B2 _3553_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_461 VGND VPWR sky130_fd_sc_hd__decap_4
X_2739_ _5292_/X _2739_/B _2740_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2900__B key_in[76] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3284__A _3284_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_645 VGND VPWR sky130_fd_sc_hd__decap_12
X_5458_ _5458_/D _2907_/A _4413_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4099__B _4098_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_133 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3306__B2 _3305_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_4409_ _4411_/A _4409_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_166 VGND VPWR sky130_fd_sc_hd__decap_6
X_5389_ _4776_/X data_out1[19] _4494_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_87_721 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3299__A1_N _3297_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_927 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_629 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_117 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3609__A2 _3607_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_960 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_971 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4843__A _4841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5233__A2_N _5258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_172 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_323 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4562__B _4557_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_654 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5231__A1 _5481_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_507 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3459__A _3459_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3237__A1_N _3257_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_520 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_721 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_907 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_564 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_743 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_406 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_586 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_236 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_235 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_664 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4742__B1 data_out1[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2810__B _2808_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_100 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_188 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3922__A _3876_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5483__RESET_B _4382_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3641__B _3640_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5412__RESET_B _4467_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_618 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_713 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_94 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3508__B1_N _3507_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_757 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_876 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_898 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_982 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_695 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3481__B1 _3465_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_643 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4025__A2 _3976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5393__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_4760_ _5490_/Q _3804_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_14_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3088__B _3088_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3784__A1 _3739_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3711_ _2717_/A _3710_/X _3741_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_159_575 VGND VPWR sky130_fd_sc_hd__fill_2
X_4691_ _2733_/C _4687_/X data_out2[8] _4688_/X _5410_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_159_597 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_3642_ _3641_/X _3642_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_247 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_718 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3536__B2 _3535_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4733__B1 data_out2[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_461 VGND VPWR sky130_fd_sc_hd__fill_2
X_3573_ _3573_/A _5516_/Q _3573_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_155_792 VGND VPWR sky130_fd_sc_hd__fill_1
X_5312_ _5297_/X _5311_/Y _5297_/X _5311_/Y _5322_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_111 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_122 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5289__A1 _3578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5289__B2 _2799_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5243_ _5233_/X _5242_/X _5233_/X _5242_/X _5243_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4928__A _4928_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_317 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3832__A _3804_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5174_ _2885_/A _5252_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_765 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_916 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3551__B key_in[31] VGND VPWR sky130_fd_sc_hd__diode_2
X_4125_ _4533_/X _4125_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_724 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5326__A1_N _5199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_4056_ _4052_/X _4055_/Y _4056_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_83_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_109 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_971 VGND VPWR sky130_fd_sc_hd__fill_1
X_3007_ _5462_/Q _3004_/X _3006_/X _3050_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_25_824 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_684 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4663__A _4518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_323 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_306 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_654 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_676 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3279__A _3213_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_389 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3224__B1 _3220_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5197__C _4679_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4958_ _4954_/Y _4958_/B _4958_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_890 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_3909_ _3062_/A _3906_/X _3908_/Y _3909_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_165_512 VGND VPWR sky130_fd_sc_hd__decap_4
X_4889_ _4886_/X _4888_/X _4889_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_20_573 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2911__A _2838_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_718 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3527__A1 _3526_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_601 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_995 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_227 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_656 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_21 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_678 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4838__A _4819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_912 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_36 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4853__B1_N _4852_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4557__B _4557_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_702 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_562 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3161__A1_N _3183_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_584 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_895 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_286 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2875__A2_N _2887_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4573__A _4573_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_738 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_749 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3189__A _3145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_827 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_996 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3215__B1 _3174_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_359 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_884 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__B1 _2973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_544 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3518__A1 data_in2[29] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_781 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5554__D _5554_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_805 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4748__A _5181_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_260 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3652__A _3579_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_794 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_540 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_670 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_746 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4483__A _4469_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_930 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3454__B1 _3438_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4914__C _4888_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_440 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3099__A _3099_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4812_ _4811_/A _4810_/X _4823_/A _4812_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_22_838 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_484 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3757__A1 _3587_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_4743_ _5481_/Q _4736_/X data_out1[2] _4737_/X _4743_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2731__A _5222_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4674_ _4674_/A _4674_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4706__B1 data_out2[14] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3509__B2 _3508_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3625_ _3618_/Y _3624_/X _3625_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__5464__D _5464_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_943 VGND VPWR sky130_fd_sc_hd__decap_3
X_3556_ _3556_/A _3555_/X _3556_/Y VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_103_604 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3390__C1 _3389_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4658__A _4525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_3487_ _3426_/X _3485_/X _3487_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_103_637 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3562__A _3562_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_125 VGND VPWR sky130_fd_sc_hd__decap_12
X_5226_ _5226_/A _5226_/B _5227_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5131__B1 _5571_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_860 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3142__C1 _3141_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_562 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_489 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1001 VGND VPWR sky130_fd_sc_hd__decap_12
X_5157_ _5154_/Y _5156_/X _5154_/Y _5156_/X _5159_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_381 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_692 VGND VPWR sky130_fd_sc_hd__decap_12
X_4108_ _4102_/Y _4105_/X _4107_/Y _4108_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_29_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_5088_ _5087_/A _5086_/Y _5096_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_779 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4237__A2 _4125_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_982 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4393__A _4390_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4039_ _4039_/A _4038_/X _4041_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3996__A1 data_in1[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_67 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_104 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_827 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_698 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_838 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_137 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_646 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1010 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4840__B _4839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_556 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2998__D _2887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_31 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3456__B _3455_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2971__A2 key_in[110] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5374__D _5374_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_773 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4568__A _4533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_326 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3472__A _3501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_979 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_860 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3191__B key_in[84] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_318 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_735 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_407 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_982 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_278 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_215 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2816__A _3778_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_440 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3987__B2 _3986_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5549__D _4545_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_771 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_473 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_782 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_635 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_821 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_523 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_820 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3647__A _5290_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_320 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_189 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5431__CLK _5430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3366__B _3362_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_352 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_363 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3371__B1_N _3370_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2962__A2 _2961_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_99 VGND VPWR sky130_fd_sc_hd__fill_2
X_3410_ _4639_/X _3404_/X _3405_/X _3406_/X _3409_/X _3410_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_4390_ _4397_/A _4390_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_171_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_902 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_602 VGND VPWR sky130_fd_sc_hd__fill_1
X_3341_ _3340_/X _3341_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_924 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4478__A _4477_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_935 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_743 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3386__B1_N _3385_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4197__B _4182_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3272_ _3268_/Y _3271_/X _3268_/Y _3271_/X _3273_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_607 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_702 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_618 VGND VPWR sky130_fd_sc_hd__fill_2
X_5011_ _4891_/A _5007_/X _5019_/B _5011_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_85_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_724 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5079__A2_N _5078_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_830 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_757 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4925__B _4924_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_513 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2726__A _2726_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_481 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5102__A _5037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4644__C _4629_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_579 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5459__D _4941_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1016 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_128 VGND VPWR sky130_fd_sc_hd__decap_3
X_2987_ _2984_/A _2984_/B _3064_/A _3065_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4726_ _4701_/A _4726_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_353 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5515__RESET_B _4344_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_898 VGND VPWR sky130_fd_sc_hd__fill_1
X_4657_ _4629_/B _4522_/A _4253_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_135_559 VGND VPWR sky130_fd_sc_hd__fill_2
X_3608_ _3608_/A _3607_/X _3608_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4588_ _3465_/A _4588_/B _4588_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_116_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3363__C1 _3362_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_710 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4388__A _4387_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3539_ _3493_/C _3539_/B _3542_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_107_34 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3292__A _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_957 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_754 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_5209_ _4635_/A _5203_/X _5204_/X _5205_/X _5208_/X _5209_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_103_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_212 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4211__A2_N _4210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_885 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_896 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_88 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_384 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3418__B1 _3403_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_473 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5454__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_977 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4570__B _4574_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_628 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_843 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_876 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_364 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5157__A1_N _5154_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3186__B _3182_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_300 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4697__A2 _4687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_784 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4298__A _4303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3633__C _5287_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_583 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_649 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3930__A _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3121__A2 key_in[114] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_852 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1010 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_576 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3409__B1 _3408_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_855 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_343 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_579 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4082__B1 _3299_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_387 VGND VPWR sky130_fd_sc_hd__decap_8
X_2910_ _2907_/X _2908_/X _2909_/Y _2910_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_90_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2691__A2_N _2690_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3890_ _3888_/X _3889_/Y _3890_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_43_292 VGND VPWR sky130_fd_sc_hd__fill_1
X_2841_ _2815_/Y _2840_/X _2815_/Y _2840_/X _2842_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_487 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3188__A2 _3186_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5560_ _5560_/D _4987_/A _4291_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2772_ _2753_/X _2771_/X _2753_/X _2771_/X _2772_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3096__B _3096_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_650 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_504 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2935__A2 key_in[109] VGND VPWR sky130_fd_sc_hd__diode_2
X_4511_ _4269_/A _4515_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_157_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_621 VGND VPWR sky130_fd_sc_hd__decap_12
X_5491_ _3836_/X _2714_/A _4373_/X _5430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_526 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_694 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4137__B2 _4136_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4442_ _4443_/A _4442_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_676 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_849 VGND VPWR sky130_fd_sc_hd__decap_12
X_4373_ _4375_/A _4373_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_421 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_966 VGND VPWR sky130_fd_sc_hd__decap_8
X_3324_ _3155_/Y _3324_/B _3324_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_59_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_977 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_988 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_573 VGND VPWR sky130_fd_sc_hd__decap_6
X_3255_ _3253_/A _3253_/B _3254_/Y _3259_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4934__A1_N _4944_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_437 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_19 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3840__A _3826_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_3186_ _3159_/B _3182_/Y _3184_/Y _3185_/Y _3186_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__4655__B _4654_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_800 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_215 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5477__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_343 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_579 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_922 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4612__A2 _4609_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_218 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3575__A1_N _5190_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4671__A _4671_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_605 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2903__B _2903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3287__A _3216_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3179__A2 _3178_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_813 VGND VPWR sky130_fd_sc_hd__fill_2
X_4709_ _5527_/Q _4699_/X data_out2[16] _4701_/X _4709_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3437__D _3436_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_846 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3734__B _3733_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3887__B1 _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_48 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5340__A3 _5337_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_732 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_99 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5007__A _5008_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_540 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_clock clkbuf_4_9_0_clock/A _5574_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_77_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_329 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4846__A _4803_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3639__B1 _3666_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3750__A _5525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_76 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_25 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4565__B _4561_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_833 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2862__A1 _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_535 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_855 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_568 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_911 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4581__A _5358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_403 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5437__RESET_B _4437_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3197__A _3125_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_84 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4906__A3 _4904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_620 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3925__A _3925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_868 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_805 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3590__A2 _3589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_849 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5562__D _4561_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_45 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3342__A2 _3340_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_936 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_81 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4756__A _4756_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3660__A _5516_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5095__A2 _5093_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3040_ _2859_/A key_in[48] _3040_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_479 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_524 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2853__A1 data_in2[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_4991_ _4992_/A _4990_/X _4991_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_63_376 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4491__A _4492_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3942_ _3941_/X _3942_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_16_292 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3819__B _3797_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2723__B _2723_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3873_ _3870_/A _3869_/X _3872_/Y _3873_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_20_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_2824_ _2968_/A key_in[42] _2824_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5543_ _5543_/D _5543_/Q _4310_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2755_ _5301_/A key_in[8] _2755_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3835__A _3835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_491 VGND VPWR sky130_fd_sc_hd__decap_12
X_5474_ _5127_/X _5116_/A _4393_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2686_ _4859_/A _2686_/B _2686_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_117_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_378 VGND VPWR sky130_fd_sc_hd__decap_4
X_4425_ _4422_/A _4425_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_890 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5472__D _5099_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3869__B1 _3866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3333__A2 _3330_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4356_ _4354_/X _4356_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1006 VGND VPWR sky130_fd_sc_hd__fill_1
X_3307_ _3299_/X _3306_/X _3299_/X _3306_/X _3318_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_424 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_724 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4666__A _4524_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_212 VGND VPWR sky130_fd_sc_hd__fill_2
X_4287_ _4289_/A _4287_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3570__A _3519_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5086__A2 _5071_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3097__A1 _3075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3238_ _3230_/X _3237_/X _3230_/X _3237_/X _3249_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_68 VGND VPWR sky130_fd_sc_hd__fill_2
X_3169_ _3169_/A _3169_/B _3170_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_54_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_855 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_814 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_151 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_836 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_23 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_549 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5530__RESET_B _4327_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_560 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_919 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_284 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_593 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_779 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_958 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_43 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_479 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_54 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3745__A _3740_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_952 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_367 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3464__B _3464_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5382__D _5382_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_860 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4576__A _4575_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_284 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3911__C _3864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2808__B _2846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_844 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_899 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_61 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2824__A _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_741 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5200__A _5200_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_713 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3260__A1 _3259_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5557__D _4554_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_757 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_222 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_256 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_266 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_621 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3655__A _3586_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_827 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2771__B1 _2762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3374__B key_in[57] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_657 VGND VPWR sky130_fd_sc_hd__decap_12
X_4210_ _4208_/X _4209_/X _4208_/X _4209_/X _4210_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_359 VGND VPWR sky130_fd_sc_hd__decap_12
X_5190_ _4798_/B _5189_/B _5211_/A _5190_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__4057__A2_N _4056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_91 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_722 VGND VPWR sky130_fd_sc_hd__decap_12
X_4141_ _4129_/Y _4159_/B _4142_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4486__A _4483_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3821__C _3820_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4072_ _4072_/A _4069_/B _4072_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_68_479 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_928 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3079__A1 _3043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2718__B _2718_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3023_ _2997_/Y _3065_/B _3023_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_343 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_899 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_674 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4028__B1 _3073_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4933__B _4932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2734__A _2733_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_4974_ _5463_/Q _4974_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5240__A2 _5209_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_3925_ _3925_/A _3924_/Y _3925_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5467__D _5035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5515__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_919 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_744 VGND VPWR sky130_fd_sc_hd__fill_2
X_3856_ data_in1[13] _3837_/X _3839_/X _3855_/Y _5492_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_165_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_407 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_2807_ _2847_/A _2847_/B _2806_/X _2846_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3003__A1 _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3787_ _3829_/A _3785_/X _3787_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_164_259 VGND VPWR sky130_fd_sc_hd__fill_2
X_5526_ _3025_/X _4707_/A _4331_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4751__A1 _4750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3554__A2 _3550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_654 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_900 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4751__B2 _4746_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2738_ _5290_/A _2737_/A _5287_/A _2943_/A _2739_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_106_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2762__B1 _2761_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3284__B _3282_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_101 VGND VPWR sky130_fd_sc_hd__fill_1
X_5457_ _4919_/X _4907_/A _4414_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_172_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_443 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_145 VGND VPWR sky130_fd_sc_hd__decap_8
X_4408_ _4411_/A _4408_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5388_ _4774_/X data_out1[18] _4495_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_733 VGND VPWR sky130_fd_sc_hd__fill_2
X_4339_ _4339_/A _4339_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4396__A _4390_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2909__A _2838_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_766 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_576 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_641 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_866 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_600 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_983 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4843__B _4842_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_994 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_471 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_538 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_869 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5020__A _5021_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5231__A2 _5229_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3459__B _3459_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3242__A1 _4718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5377__D _4752_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4135__A1_N _4133_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_733 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_576 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_766 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_737 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_247 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4742__A1 _3583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4742__B2 _4737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2810__C _2809_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_613 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2753__B1 _2801_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_793 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3922__B _3922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_690 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2819__A _2819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_381 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_906 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_clock clkbuf_2_2_0_clock/X clkbuf_3_5_0_clock/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_19_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_896 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_961 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5452__RESET_B _4420_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_888 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_365 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3481__B2 _3480_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5538__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_847 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_3710_ _3702_/Y _3709_/X _3710_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__3784__A2 _3783_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4690_ _5518_/Q _4687_/X data_out2[7] _4688_/X _4690_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_14_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_92 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_3641_ _3641_/A _3640_/X _3641_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_128_941 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3385__A _4728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_708 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4733__A1 _5539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3572_ _5516_/Q _3572_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4733__B2 _4726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_996 VGND VPWR sky130_fd_sc_hd__fill_2
X_5311_ _5306_/Y _5308_/X _5310_/Y _5311_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_142_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_977 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5289__A2 _5288_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_808 VGND VPWR sky130_fd_sc_hd__fill_2
X_5242_ _5239_/X _5241_/B _5241_/X _5242_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_130_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_796 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4928__B _4927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_178 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3832__B _3832_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_329 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2729__A _2852_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5173_ _5355_/A _2885_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_60_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_841 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5105__A _5104_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_608 VGND VPWR sky130_fd_sc_hd__fill_2
X_4124_ data_in1[24] _3976_/X _4091_/X _4123_/Y _5503_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_84_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4249__B1 _4248_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_118 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_4055_ _4030_/Y _4053_/Y _4054_/Y _4055_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4944__A _4944_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_630 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_3006_ _3052_/A _3052_/B _3006_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_83_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4663__B _4521_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_633 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_308 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_132 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_319 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_143 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3279__B _3244_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_688 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3224__A1 _4638_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4957_ _4554_/A _4956_/X _4554_/A _4956_/X _4958_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3224__B2 _3223_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3908_ _3908_/A _3908_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4888_ _4865_/X _4877_/X _4866_/X _4875_/X _4887_/Y _4888_/X VGND VPWR sky130_fd_sc_hd__o32a_4
XFILLER_138_727 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2983__B1 _2998_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3839_ _3839_/A _3812_/B _3875_/A _3839_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__2911__B _2865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_941 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3527__A2 _3526_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_922 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_613 VGND VPWR sky130_fd_sc_hd__decap_12
X_5509_ _5509_/D _3368_/A _4351_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4838__B _4838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_924 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_48 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5015__A _4975_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_852 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_928 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_574 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4854__A _4840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2839__B1_N _2838_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_769 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_825 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4573__B _4561_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3189__B key_in[52] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_85 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_463 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3215__A1 data_in2[20] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_705 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__A1 _4870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__B2 _4930_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_738 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_524 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_51 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2974__B1 _2973_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_226 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_40 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3518__A2 _3391_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_730 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_741 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_977 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4012__A1_N _3999_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_762 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_487 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_947 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3652__B _3650_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5570__D _5570_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_585 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1001 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_994 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3454__B2 _3464_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3099__B _3099_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4811_ _4811_/A _4810_/X _4823_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_61_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_891 VGND VPWR sky130_fd_sc_hd__decap_6
X_4742_ _3583_/C _4736_/X data_out1[1] _4737_/X _5371_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3757__A2 _3737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_861 VGND VPWR sky130_fd_sc_hd__decap_3
X_4673_ _4672_/X _4674_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_30_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_708 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4706__A1 _2984_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3624_ _3624_/A _3623_/X _3624_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__4706__B2 _4701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4004__A _3957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_590 VGND VPWR sky130_fd_sc_hd__decap_12
X_3555_ _5164_/Y _3554_/Y _5164_/Y _3554_/Y _3555_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_432 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4939__A _4938_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3843__A _3721_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_817 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_914 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5232__A2_N _5361_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3390__B1 _3364_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_999 VGND VPWR sky130_fd_sc_hd__decap_8
X_3486_ _3429_/B _3485_/X _3488_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_142_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4658__B _4586_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3562__B _3562_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_5225_ _5513_/Q _3603_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_103_649 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_435 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5480__D _3598_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5131__B2 _5130_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3142__B1 _3103_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5374__RESET_B _4512_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_405 VGND VPWR sky130_fd_sc_hd__fill_2
X_5156_ _4573_/A _5155_/X _4573_/A _5155_/X _5156_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3866__A1_N _2980_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_4107_ _4106_/X _4107_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_110_170 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4674__A _4674_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5087_ _5087_/A _5086_/Y _5087_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_84_577 VGND VPWR sky130_fd_sc_hd__decap_3
X_4038_ _4778_/X _4036_/X _4037_/X _4038_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_25_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3996__A2 _3976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_290 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_17 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_806 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_305 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_658 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2922__A _2849_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_343 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_376 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2708__B1 _5303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_410 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4849__A _5547_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_559 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_977 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3381__B1 _3341_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_593 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3472__B key_in[92] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5383__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5390__D _4777_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_446 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_872 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_371 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4881__B1 _4871_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_747 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4584__A _4521_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_514 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_62 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_599 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4633__B1 _4800_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_482 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_666 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_50 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2832__A _2832_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4936__A1 _4642_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_72 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_833 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3647__B _3646_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2947__B1 _2939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_894 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5565__D _4564_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_843 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_320 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_888 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_376 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_538 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_869 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3663__A _3662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_3340_ _5076_/A _3340_/B _3340_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_113_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_614 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_958 VGND VPWR sky130_fd_sc_hd__decap_8
X_3271_ _3270_/X _3271_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_809 VGND VPWR sky130_fd_sc_hd__decap_12
X_5010_ _5009_/X _5019_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_23_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_883 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_894 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_371 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4494__A _4492_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A clkbuf_2_2_0_clock/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_39_769 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_341 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_536 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5102__B _5101_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_953 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_441 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_625 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3838__A _4537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_800 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_669 VGND VPWR sky130_fd_sc_hd__decap_12
X_2986_ _2986_/A _3064_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_148_811 VGND VPWR sky130_fd_sc_hd__decap_12
X_4725_ _4699_/A _4725_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5475__D _5142_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_4656_ _4655_/X _4656_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_376 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2874__A2_N _2873_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3607_ _3601_/Y _3606_/X _3601_/Y _3606_/X _3607_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_730 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4669__A _4631_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4587_ _4518_/X _4629_/B _4578_/A _4586_/X _4588_/B VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3573__A _3573_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_379 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3363__B1 _3316_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_560 VGND VPWR sky130_fd_sc_hd__fill_2
X_3538_ _3521_/X _3537_/X _3521_/X _3537_/X _3543_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5555__RESET_B _4296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_582 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_733 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3292__B key_in[23] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_947 VGND VPWR sky130_fd_sc_hd__decap_4
X_3469_ _3469_/A _3468_/X _3469_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_89_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_5208_ _5234_/A key_in[97] _5303_/A _5208_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_88_179 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_680 VGND VPWR sky130_fd_sc_hd__decap_12
X_5139_ _5133_/Y _5140_/B _5139_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3418__B2 _3417_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_238 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_953 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_98 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3748__A _3765_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_1008 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_4_0_clock clkbuf_4_5_0_clock/A _5530_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__5040__B1 _5564_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_855 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5385__D _4768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3186__C _3184_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3758__A1_N _3756_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_398 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_741 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4579__A _4579_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_508 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_345 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_378 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_52 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3106__B1 _2999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3930__B _3925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2827__A _2898_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_864 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5203__A _5203_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_363 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3409__A1 _3499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_322 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_964 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4082__B2 _4081_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_591 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3658__A _3681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_619 VGND VPWR sky130_fd_sc_hd__fill_2
X_2840_ _2840_/A _2839_/X _2840_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_148_107 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5031__B1 _5017_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_129 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _2762_/Y _2770_/Y _2762_/Y _2770_/Y _2771_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_691 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_803 VGND VPWR sky130_fd_sc_hd__fill_2
X_4510_ _4504_/X _4510_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_156_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_662 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3593__B1 _3587_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5490_ _3810_/X _5490_/Q _4374_/X _5430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_157_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_538 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_633 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_195 VGND VPWR sky130_fd_sc_hd__decap_3
X_4441_ _4443_/A _4441_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4489__A _4483_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3393__A _3519_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_912 VGND VPWR sky130_fd_sc_hd__decap_3
X_4372_ _4375_/A _4372_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_153_891 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_582 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_3323_ _3180_/A _3322_/A _3010_/A _3495_/B _3324_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_98_433 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_777 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_265 VGND VPWR sky130_fd_sc_hd__decap_8
X_3254_ _3305_/A _3254_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_101_939 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3648__A1 _5290_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5202__A1_N _5181_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4845__B1 _4836_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3840__B _3833_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_842 VGND VPWR sky130_fd_sc_hd__decap_4
X_3185_ _3112_/X _3185_/B _3185_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2737__A _2737_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_190 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5113__A _5113_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4952__A _4918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_761 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4671__B _4656_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_794 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3568__A _4664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_591 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_956 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3557__A2_N _3556_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_967 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_416 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5022__B1 _5017_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_617 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3287__B _3143_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2969_ _2934_/A key_in[14] _2969_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4708_ _3020_/A _4699_/X data_out2[15] _4701_/X _4708_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_136_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_858 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4399__A _4402_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4639_ _4638_/X _4639_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_151_806 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_817 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_327 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3887__A1 _3682_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3887__B2 _3175_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_849 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5007__B _5006_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_744 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_232 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5089__B1 _5076_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_563 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3639__A1 _5284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_609 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5023__A _5023_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5421__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_300 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2862__A2 key_in[107] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_86 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_388 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_400 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_591 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5571__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3197__B _3197_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_641 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_961 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_803 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_96 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3575__B1 _5190_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5477__RESET_B _4389_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_847 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_110 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3925__B _3924_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5406__RESET_B _4474_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_120 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3327__B1 _3326_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_676 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_582 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_861 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_606 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_959 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3660__B _3659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5016__A2_N _5015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_834 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_620 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2853__A2 _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4772__A _2889_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4990_ _4978_/Y _4983_/B _4990_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_90_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_539 VGND VPWR sky130_fd_sc_hd__fill_2
X_3941_ _3938_/X _3940_/X _3938_/X _3940_/X _3941_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_731 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3388__A _3388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_416 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_3872_ _3871_/X _3872_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_31_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5004__B1 _4978_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_797 VGND VPWR sky130_fd_sc_hd__decap_12
X_2823_ _2822_/A _2821_/X _2822_/X _2840_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_20_959 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3566__B1 data_in2[31] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_803 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_814 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_2754_ _5300_/A key_in[40] _2754_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5542_ _3567_/Y _5542_/Q _4312_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_118_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_982 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_493 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4210__A2_N _4209_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_644 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3835__B _3833_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_858 VGND VPWR sky130_fd_sc_hd__decap_4
X_5473_ _5115_/X _5473_/Q _4394_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_133_806 VGND VPWR sky130_fd_sc_hd__fill_2
X_2685_ _4636_/A _5366_/X _5367_/X _5368_/X _5369_/X _2686_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_144_154 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5108__A _5087_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4424_ _4422_/A _4424_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_699 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3869__B2 _3868_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_349 VGND VPWR sky130_fd_sc_hd__decap_4
X_4355_ _4354_/X _4355_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_764 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4947__A _4943_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_19 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3851__A _3875_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3306_ _3304_/X _3305_/X _3304_/X _3305_/X _3306_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_403 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_574 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5444__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4286_ _4289_/A _4286_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4666__B _4629_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_436 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3570__B _3570_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5086__A3 _5058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_758 VGND VPWR sky130_fd_sc_hd__fill_2
X_3237_ _3257_/B _3236_/X _3257_/B _3236_/X _3237_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_650 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3481__A2_N _3480_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3097__A2 _3095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_25 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_514 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_300 VGND VPWR sky130_fd_sc_hd__decap_6
X_3168_ _3169_/A _3169_/B _3170_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_67_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_536 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5156__A1_N _4573_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_845 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_642 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3099_ _3099_/A _3099_/B _3099_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5243__B1 _5233_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_366 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_539 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_703 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_725 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_904 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_736 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_202 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_274 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_425 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_961 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_22 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3557__B1 _3548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2930__A _2930_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5570__RESET_B _4279_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3745__B _3742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_625 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_880 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4857__A _4857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_872 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3761__A _3749_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2690__A2_N _2689_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_414 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_447 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_801 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_108 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_837 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_697 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_314 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_848 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2824__B key_in[42] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3796__B1 _5518_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_753 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_550 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3260__A2 _3258_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3001__A _2790_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_274 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_clock clkbuf_2_0_0_clock/X clkbuf_4_3_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_9_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2840__A _2840_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_931 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_493 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_953 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_964 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5573__D _4573_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2771__B2 _2770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_934 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5467__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_349 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_669 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4767__A _5494_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_904 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3671__A _3671_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4140_ _4129_/Y _4159_/B _4142_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3720__B1 _3681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_948 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_734 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_544 VGND VPWR sky130_fd_sc_hd__decap_12
X_4071_ _4026_/A _3950_/B _4784_/X _4071_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3079__A2 key_in[113] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_577 VGND VPWR sky130_fd_sc_hd__decap_3
X_3022_ _2997_/Y _3065_/B _3022_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_49_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4028__A1 _3075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_984 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4028__B2 _3394_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_4973_ _4870_/X _4971_/X _4972_/Y _5462_/Q _4930_/X _5462_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__5399__RESET_B _4482_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3924_ _3895_/X _3920_/Y _3922_/Y _3923_/Y _3924_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__4984__C1 _4983_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4007__A _3959_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_892 VGND VPWR sky130_fd_sc_hd__decap_12
X_3855_ _3835_/A _3853_/Y _3854_/X _3855_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_20_756 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2750__A _2742_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2806_ _2847_/A _2847_/B _2806_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_164_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_3786_ _3829_/A _3785_/X _3786_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3003__A2 key_in[111] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_953 VGND VPWR sky130_fd_sc_hd__fill_1
X_5525_ _5525_/D _5525_/Q _4332_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4751__A2 _4745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3554__A3 _3551_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5483__D _3653_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2737_ _2737_/A _2943_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_986 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2762__A1 _4882_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_934 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_176 VGND VPWR sky130_fd_sc_hd__fill_2
X_5456_ _4906_/Y _5456_/Q _4415_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_956 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5161__C1 _5160_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4407_ _4411_/A _4407_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4677__A _4677_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_550 VGND VPWR sky130_fd_sc_hd__decap_3
X_5387_ _4773_/X data_out1[17] _4496_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3581__A _5222_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_872 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_583 VGND VPWR sky130_fd_sc_hd__fill_2
X_4338_ _4339_/A _4338_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2909__B _2865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_522 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_458 VGND VPWR sky130_fd_sc_hd__fill_1
X_4269_ _4269_/A _4271_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_47_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_801 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_588 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_940 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2925__A _2925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2721__A1_N _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_878 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_506 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_815 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5216__B1 _4679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5301__A _5301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_16 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_848 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_859 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5020__B _5019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_870 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3242__A2 _3280_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_572 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_881 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_65 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_892 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_233 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_705 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_739 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_920 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_964 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5393__D _4785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3373__A2_N _3372_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4742__A2 _4736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_259 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_912 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_219 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2753__A1 _2742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_410 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_944 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_809 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4587__A _4518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_466 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_977 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3491__A _3317_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_62 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2819__B _2819_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_95 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_918 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_704 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_823 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_642 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2835__A _4900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3941__A2_N _3940_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_973 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_83 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5211__A _5211_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_377 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_859 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5568__D _4567_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_196 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5492__RESET_B _4372_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5421__RESET_B _4457_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_717 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3666__A _3666_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3640_ _5253_/Y _2735_/X _3624_/A _3621_/X _3640_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_146_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3385__B _3385_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3571_ _3676_/A _3579_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_901 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4733__A2 _4725_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_5310_ _5309_/X _5310_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3941__B1 _3938_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_422 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_793 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_5241_ _5239_/X _5241_/B _5241_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_455 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4497__A _4269_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_989 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_308 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_499 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3832__C _3830_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5172_ _5172_/A _5355_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_520 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2729__B _2727_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_745 VGND VPWR sky130_fd_sc_hd__decap_12
X_4123_ _4092_/X _4123_/B _4123_/C _4123_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_111_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_564 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4249__A1 _4246_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_288 VGND VPWR sky130_fd_sc_hd__fill_1
X_4054_ _4003_/X _4031_/X _4008_/Y _4054_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_110_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4944__B _4932_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3005_ _3004_/X _3052_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_37_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_269 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2745__A _2744_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5121__A _5121_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4663__C _4523_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_848 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5509__RESET_B _4351_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_196 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5478__D _5171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_291 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4960__A _4947_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_829 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_4956_ _4921_/X _4955_/X _4956_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3224__A2 _3218_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_188 VGND VPWR sky130_fd_sc_hd__fill_2
X_3907_ _3062_/A _3906_/X _3908_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_4887_ _4864_/Y _4887_/B _4887_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3576__A _3575_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_739 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2983__B2 _2982_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3838_ _4537_/X _3839_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_165_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2911__C _2834_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_953 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_761 VGND VPWR sky130_fd_sc_hd__fill_2
X_3769_ _2842_/A _3769_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_452 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_934 VGND VPWR sky130_fd_sc_hd__decap_12
X_5508_ _5508_/D _3322_/A _4352_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_106_625 VGND VPWR sky130_fd_sc_hd__decap_12
X_5439_ _4592_/X _4589_/A _4435_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_121_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4200__A _4178_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_680 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3696__C1 _3695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_542 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5015__B _5014_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_864 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_299 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4854__B _4844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_623 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_943 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5388__D _4774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_111 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_280 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_656 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_667 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4870__A _4857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_987 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3215__A2 _3172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_328 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_531 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__A2 _4961_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__A _3429_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_897 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_374 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_728 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2974__A1 _2973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_385 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_575 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_524 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_249 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4176__B1 _3452_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_989 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_774 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5206__A _5203_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_317 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_499 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4110__A _4109_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3652__C _3651_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_907 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5505__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_417 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_597 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_940 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_111 VGND VPWR sky130_fd_sc_hd__decap_8
X_4810_ _4837_/B _4810_/B _4810_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__4780__A _3085_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_987 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_497 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_330 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_380 VGND VPWR sky130_fd_sc_hd__decap_12
X_4741_ _5480_/Q _3583_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3396__A _3231_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_525 VGND VPWR sky130_fd_sc_hd__decap_12
X_4672_ _4671_/X _4672_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4706__A2 _4699_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3623_ _5272_/Y _3622_/X _5272_/Y _3622_/X _3623_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_750 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_761 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4004__B _3982_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_912 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_271 VGND VPWR sky130_fd_sc_hd__fill_2
X_3554_ _4640_/X _3550_/X _3551_/X _3552_/X _3553_/X _3554_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XANTENNA__4939__B _4937_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_753 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3843__B _3841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3390__A1 data_in2[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_444 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_455 VGND VPWR sky130_fd_sc_hd__fill_2
X_3485_ _3431_/A _3459_/B _3485_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_786 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_477 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5116__A _5116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4658__C _4519_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_328 VGND VPWR sky130_fd_sc_hd__decap_8
X_5224_ _5252_/A _5252_/B _5513_/Q _5224_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__4020__A _4020_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_296 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_840 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3142__A1 data_in2[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_149 VGND VPWR sky130_fd_sc_hd__decap_4
X_5155_ _4572_/A _5052_/A _5144_/X _5155_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4955__A _4553_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_575 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_737 VGND VPWR sky130_fd_sc_hd__fill_2
X_4106_ _4102_/Y _4105_/X _4106_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_5086_ _5059_/A _5071_/Y _5058_/X _5084_/Y _5085_/X _5086_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_110_182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_247 VGND VPWR sky130_fd_sc_hd__fill_1
X_4037_ _4778_/X _4036_/X _4037_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_71_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_36 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_280 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_656 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_29 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_615 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_149 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2922__B _2921_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4939_ _4938_/A _4937_/X _4949_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_895 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4158__B1 _4157_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_517 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_761 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2708__A1 _5299_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_388 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_783 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_77 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4849__B _4838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_549 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_956 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3381__A1 _3342_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5528__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_989 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_797 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_425 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_clock clkbuf_4_1_0_clock/A _5498_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_153_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_501 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_361 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_76 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4881__A1 _4870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4881__B2 _4815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_940 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_450 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4633__A1 _3529_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_472 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4633__B2 _4631_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_228 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_239 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_420 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_188 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_659 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4936__A2 _4934_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_503 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_851 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2947__B2 _2946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_845 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_13 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_310 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_332 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_580 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_414 VGND VPWR sky130_fd_sc_hd__fill_2
X_3270_ _3227_/A _3269_/Y _3270_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_3_593 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4775__A _2959_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_854 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_707 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_461 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_272 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2823__B1_N _2822_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_659 VGND VPWR sky130_fd_sc_hd__decap_3
X_2985_ _2984_/X _2986_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_823 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2938__A1 _4943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_171 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4015__A _3972_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4724_ _5535_/Q _3316_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_159_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_322 VGND VPWR sky130_fd_sc_hd__fill_2
X_4655_ _4809_/B _4654_/Y _4655_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_388 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3854__A _3840_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_539 VGND VPWR sky130_fd_sc_hd__fill_2
X_3606_ _3619_/A _3605_/X _3619_/A _3605_/X _3606_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_347 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4669__B _4662_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4586_ _4524_/A _4586_/B _4586_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_742 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3573__B _5516_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3363__A1 data_in2[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5491__D _3836_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3537_ _3522_/X _3536_/X _3522_/X _3536_/X _3537_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_594 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_648 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_659 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_436 VGND VPWR sky130_fd_sc_hd__fill_2
X_3468_ _3108_/Y _3251_/Y _3441_/X _3468_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_131_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_244 VGND VPWR sky130_fd_sc_hd__fill_1
X_5207_ _5207_/A _5303_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_350 VGND VPWR sky130_fd_sc_hd__decap_12
X_3399_ _3231_/Y _3398_/X _3399_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_692 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5524__RESET_B _4334_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5138_ _5138_/A _5138_/B _5136_/Y _5137_/Y _5140_/B VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2874__B1 _3801_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_5069_ _5068_/X _5084_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2933__A _2934_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_773 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_615 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4011__A1_N _3200_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_637 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3748__B _3679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_648 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_467 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5040__B2 _5039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3186__D _3185_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_377 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_814 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_314 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_76 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_847 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_357 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_103 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_211 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3106__A1 _3060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4989__B1_N _4988_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_552 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4595__A _5441_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_117 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_331 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_707 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4912__B1_N _4911_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_876 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5203__B key_in[33] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_824 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3409__A2 key_in[122] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_442 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3939__A _3794_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3850__A1_N _3847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_987 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_773 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2843__A _2842_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_434 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3658__B _3680_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_979 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5576__D _5576_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5031__A1 _5001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5031__B2 _5017_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_620 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_631 VGND VPWR sky130_fd_sc_hd__decap_4
X_2770_ _2770_/A _2770_/B _2768_/X _2769_/Y _2770_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2949__A2_N _2948_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4790__B1 data_out1[26] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3593__B2 _3592_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_837 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3674__A _3674_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4440_ _4419_/A _4443_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_172_645 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_195 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3393__B _3364_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_818 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_561 VGND VPWR sky130_fd_sc_hd__decap_4
X_4371_ _4375_/A _4371_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_701 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_3322_ _3322_/A _3495_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_4_891 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_445 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_478 VGND VPWR sky130_fd_sc_hd__decap_12
X_3253_ _3253_/A _3253_/B _3305_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_789 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4845__A1 _4802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3648__A2 _3646_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_428 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3803__A1_N _3794_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4845__B2 _4815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_832 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1011 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_534 VGND VPWR sky130_fd_sc_hd__fill_2
X_3184_ _3115_/B _3185_/B _3184_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_39_556 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5113__B _5111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_898 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3506__B1_N _3477_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_846 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4952__B _4950_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_367 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_570 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3281__B1 _3241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4671__C _4659_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_890 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_732 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5486__D _3718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5022__A1 _4896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5373__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_776 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5022__B2 _4806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3287__C _3287_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_631 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_629 VGND VPWR sky130_fd_sc_hd__fill_1
X_2968_ _2968_/A key_in[46] _2968_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_148_642 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2777__B1_N _2776_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4707_ _4707_/A _3020_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_163_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3584__A _4524_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2899_ _2790_/A key_in[12] _2899_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_163_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_174 VGND VPWR sky130_fd_sc_hd__decap_4
X_4638_ _4637_/X _4638_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4569_ _5569_/Q _4574_/B _5569_/D VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3887__A2 _3175_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5089__A1 _4870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5089__B2 _4930_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3639__A2 _3638_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_846 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_194 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3759__A _3759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3272__B1 _3268_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_710 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_743 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_31 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_754 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5396__D _4790_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_467 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3197__C _3129_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3575__B2 _3574_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3327__A1 _3155_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3602__A2_N _3589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_870 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_520 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5446__RESET_B _4427_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_715 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2838__A _2838_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_748 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_662 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_813 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_684 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2873__A2_N _2872_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_751 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5396__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_762 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_367 VGND VPWR sky130_fd_sc_hd__decap_3
X_3940_ _3939_/X _3904_/X _3916_/X _3940_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_44_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_743 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3388__B _3388_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3871_ _3870_/X _3871_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5004__A1 _4985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_2822_ _2822_/A _2821_/X _2822_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_31_275 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_297 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3566__A1 _5197_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5541_ _3546_/X _5541_/Q _4313_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3566__B2 _4546_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2753_ _2742_/X _2749_/Y _2801_/B _2753_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_145_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_471 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3835__C _3834_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5472_ _5099_/Y _5472_/Q _4395_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4423_ _4422_/A _4423_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5108__B _5098_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_497 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_188 VGND VPWR sky130_fd_sc_hd__decap_12
X_4354_ _4340_/A _4354_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4947__B _4946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3851__B _3850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_916 VGND VPWR sky130_fd_sc_hd__decap_6
X_3305_ _3305_/A _3305_/B _3305_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_140_361 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2748__A _5332_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_798 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_4285_ _4289_/A _4285_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_949 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_586 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5124__A _5124_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4666__C _4518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_597 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3570__C _3577_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3236_ _3236_/A _3187_/X _3236_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_86_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2829__B1 _2828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_247 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_802 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_813 VGND VPWR sky130_fd_sc_hd__decap_12
X_3167_ _3143_/C _3166_/B _3166_/X _3169_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_95_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_194 VGND VPWR sky130_fd_sc_hd__decap_12
X_3098_ _3099_/A _3099_/B _3098_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_507 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3579__A _3579_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5243__B2 _5242_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_710 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_592 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_69 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_776 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_916 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_748 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_225 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_23 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_437 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3557__B2 _3556_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2930__B _2925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_612 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_494 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4203__A _4092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_965 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_78 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_464 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4857__B _4855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_669 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3761__B _3782_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_884 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5034__A _5034_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_813 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4873__A _4873_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_97 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4977__A2_N _4976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_632 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3489__A _3489_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3796__A1 _2723_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_220 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3796__B2 _3062_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3001__B key_in[15] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_286 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_595 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_770 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2840__B _2839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_781 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_931 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4113__A _4068_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_964 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_975 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_166 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_997 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5216__A1_N _4679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3952__A _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_328 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_916 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3671__B _3670_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3720__A1 _3701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_437 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_394 VGND VPWR sky130_fd_sc_hd__decap_3
X_4070_ data_in1[22] _3976_/X _4043_/X _4069_/Y _4070_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_68_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_556 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_651 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_960 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_802 VGND VPWR sky130_fd_sc_hd__decap_12
X_3021_ _3021_/A _3020_/Y _3065_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_48_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_589 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4175__B1_N _4174_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4028__A2 _5537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3399__A _3231_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_849 VGND VPWR sky130_fd_sc_hd__decap_4
X_4972_ _4971_/A _4970_/X _4972_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_3923_ _3874_/X _3922_/B _3923_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4984__B1 _4942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_540 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4007__B _4007_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2995__C1 _2994_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_882 VGND VPWR sky130_fd_sc_hd__decap_3
X_3854_ _3840_/Y _3852_/X _3854_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2805_ _2814_/D _2804_/X _2814_/D _2804_/X _2847_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__2750__B _2749_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1004 VGND VPWR sky130_fd_sc_hd__decap_3
X_3785_ _3831_/A _3785_/B _3785_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_164_239 VGND VPWR sky130_fd_sc_hd__decap_4
X_5524_ _5524_/D _5524_/Q _4334_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4023__A _4014_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2736_ _2702_/X _2722_/B _5358_/A _2736_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3509__A2_N _3508_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5411__CLK _5402_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_667 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_998 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2762__A2 _2759_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_261 VGND VPWR sky130_fd_sc_hd__decap_12
X_5455_ _5455_/D _4882_/A _4416_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_626 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4958__A _4954_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_497 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3862__A _3817_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_968 VGND VPWR sky130_fd_sc_hd__decap_8
X_4406_ _4411_/A _4406_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5161__B1 _4542_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5386_ _4771_/X data_out1[16] _4498_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_1005 VGND VPWR sky130_fd_sc_hd__fill_2
X_4337_ _4339_/A _4337_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5561__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2909__C _2836_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_534 VGND VPWR sky130_fd_sc_hd__decap_12
X_4268_ _4267_/Y _4269_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_28_813 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_150 VGND VPWR sky130_fd_sc_hd__fill_2
X_3219_ _3148_/A key_in[21] _3219_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3475__B1 _5128_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4199_ _4159_/X _4198_/B _4200_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_83_952 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_963 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2925__B _2924_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5216__B2 _5215_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_367 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5301__B key_in[4] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3102__A _5355_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_501 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_562 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_584 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_77 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4727__B1 data_out2[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_770 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_728 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_227 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2753__A2 _2749_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4868__A _4865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3772__A _3769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_497 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5152__B1 _5132_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_967 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4587__B _4629_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_851 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3491__B _3491_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_862 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_835 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_846 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_51 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2835__B _2794_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_805 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5211__B _5210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_687 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_698 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3012__A _3012_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_348 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_871 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3947__A _3835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_573 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2851__A _2850_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5434__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3666__B _3666_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3480__A2_N _3479_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_239 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_291 VGND VPWR sky130_fd_sc_hd__decap_3
X_3570_ _3519_/A _3570_/B _3577_/A _3570_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5461__RESET_B _4409_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_762 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_913 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4239__A2_N _3556_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_250 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4778__A _3030_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3941__B2 _3940_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_721 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_260 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3682__A _5522_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_968 VGND VPWR sky130_fd_sc_hd__decap_8
X_5240_ _4811_/A _5209_/Y _5211_/X _5241_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_5_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_670 VGND VPWR sky130_fd_sc_hd__fill_1
X_5171_ _5478_/Q _4995_/X _4542_/B _5170_/Y _5171_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3832__D _3831_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2729__C _2728_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_4122_ _4112_/X _4120_/Y _4123_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_69_757 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4249__A2 _4247_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_576 VGND VPWR sky130_fd_sc_hd__decap_4
X_4053_ _4002_/X _4029_/X _4053_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_83_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_481 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_790 VGND VPWR sky130_fd_sc_hd__decap_3
X_3004_ _4637_/A _3000_/X _3001_/X _3002_/X _3003_/X _3004_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_65_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_676 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4663__D _4586_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_911 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5121__B _5119_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_996 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4018__A _3966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_101 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_27 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4957__B1 _4554_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4955_ _4553_/A _4944_/X _4955_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4960__B _4950_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3857__A _3839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3224__A3 _3219_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2761__A _2761_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3906_ _2918_/A _3905_/A _5523_/Q _3905_/Y _3906_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__5549__RESET_B _4303_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4886_ _4885_/A _4884_/X _4885_/Y _4886_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_60_690 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4709__B1 data_out2[16] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5494__D _5494_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3837_ _4533_/X _3837_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_165_526 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3448__A2_N _3447_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2911__D _2770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3768_ _3681_/A _3767_/X _3768_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_119_965 VGND VPWR sky130_fd_sc_hd__decap_6
X_5507_ _4204_/X _3300_/A _4353_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4688__A _4677_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_710 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_208 VGND VPWR sky130_fd_sc_hd__fill_2
X_2719_ _2719_/A _5364_/X _2719_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3699_ _3765_/A _3679_/B _5229_/A _3699_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_106_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_648 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_46 VGND VPWR sky130_fd_sc_hd__decap_4
X_5438_ _4643_/Y _4635_/A _4436_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_979 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_24 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_57 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_670 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_286 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_68 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4200__B _4196_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5369_ _5300_/A key_in[102] _2828_/A _5369_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3696__B1 _3679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_256 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_876 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_407 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3448__B1 _5116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_10 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5457__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1007 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_966 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_871 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__A _3701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3620__B1 _3619_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__A3 _4962_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_543 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__B _3485_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_515 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2974__A2 _2972_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_587 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4176__B2 _4175_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_329 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_990 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_50 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_204 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_738 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2846__A _2778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3439__B1 _3108_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_226 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_749 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5222__A _5222_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_237 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_120 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_665 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5579__D _4264_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_432 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_4740_ _3577_/A _4736_/X data_out1[0] _4737_/X _4740_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_14_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_4671_ _4671_/A _4656_/X _4659_/Y _4670_/X _4671_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_147_537 VGND VPWR sky130_fd_sc_hd__decap_12
X_3622_ _5514_/Q _2733_/C _3621_/X _3622_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3914__A1 _3909_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3553_ _3528_/A key_in[127] _3408_/X _3553_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_116_935 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2720__A1_N _2744_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_220 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4301__A _4303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3390__A2 _3172_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3484_ _3484_/A _3457_/B _3488_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_131_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_5223_ _5223_/A _5252_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_798 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4658__D _4253_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4020__B _4018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3142__A2 _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_852 VGND VPWR sky130_fd_sc_hd__fill_2
X_5154_ _5477_/Q _5154_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_651 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4955__B _4944_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_513 VGND VPWR sky130_fd_sc_hd__fill_2
X_4105_ _4051_/Y _4103_/Y _4078_/Y _4104_/Y _4105_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_56_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2756__A _5301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_684 VGND VPWR sky130_fd_sc_hd__fill_2
X_5085_ _5072_/A _5085_/B _5085_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5132__A _5132_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_194 VGND VPWR sky130_fd_sc_hd__decap_12
X_4036_ _4034_/X _4035_/X _4034_/X _4035_/X _4036_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_451 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_900 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5489__D _3789_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_782 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4971__A _4971_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_635 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3850__B1 _3847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5365__B1_N _5364_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_977 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_465 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_167 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_785 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3587__A _3575_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5383__RESET_B _4501_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4938_ _4938_/A _4937_/X _4938_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3602__B1 _3573_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_830 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_835 VGND VPWR sky130_fd_sc_hd__decap_4
X_4869_ _4802_/X _4867_/Y _4868_/X _4859_/A _4815_/X _4869_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4158__A1 _3396_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_751 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_529 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2708__A2 key_in[103] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_250 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_34 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5307__A _4827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_89 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_220 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5107__B1 _5124_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_968 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_294 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3381__A2 _3346_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_938 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_329 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_415 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3669__B1 _3665_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_66 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4881__A2 _4879_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_161 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2892__A1 _2714_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5042__A _5041_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_719 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5399__D _5399_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_613 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4633__A2 _4631_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_730 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3841__B1 _2847_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_432 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_741 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_999 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_651 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_684 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_863 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_312 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_526 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_537 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5346__B1 _5335_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_384 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_344 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_272 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_399 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_294 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5217__A _5192_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4121__A _4112_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_735 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3960__A _3073_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_768 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_502 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_760 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4085__B1 _4115_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5282__C1 _5281_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_473 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4791__A _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_421 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_741 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_966 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_925 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_958 VGND VPWR sky130_fd_sc_hd__decap_12
X_2984_ _2984_/A _2984_/B _2984_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4723_ _3287_/C _4712_/X data_out2[23] _4713_/X _5425_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2938__A2 _2936_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4015__B _4015_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4654_ _4525_/X _4586_/B _4519_/X _4666_/D _4654_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_147_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_827 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_838 VGND VPWR sky130_fd_sc_hd__decap_4
X_3605_ _5242_/X _3604_/Y _5242_/X _3604_/Y _3605_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3854__B _3852_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_4585_ _4650_/B _4586_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_162_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4669__C _3676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_359 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3418__A1_N _3403_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_754 VGND VPWR sky130_fd_sc_hd__decap_8
X_3536_ _3527_/X _3535_/X _3527_/X _3535_/X _3536_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4031__A _4029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3363__A2 _3172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_702 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_404 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_724 VGND VPWR sky130_fd_sc_hd__decap_4
X_3467_ _4786_/X _3300_/A _3466_/X _3469_/A VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__4966__A _4921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3870__A _3870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_297 VGND VPWR sky130_fd_sc_hd__decap_8
X_5206_ _5203_/A _5234_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_779 VGND VPWR sky130_fd_sc_hd__decap_12
X_3398_ _3253_/A _5510_/Q _4043_/C _3397_/Y _3398_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_97_660 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_971 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_362 VGND VPWR sky130_fd_sc_hd__decap_4
X_5137_ _5108_/X _5137_/B _5086_/Y _5137_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_112_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_395 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_321 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2874__B2 _2873_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_708 VGND VPWR sky130_fd_sc_hd__decap_8
X_5068_ _5068_/A _5067_/X _5068_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_888 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2689__A1_N _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4076__B1 _3143_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_771 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_922 VGND VPWR sky130_fd_sc_hd__decap_12
X_4019_ _3970_/Y _4019_/B _4019_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_84_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5564__RESET_B _4286_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_730 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3823__B1 _2914_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_903 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_988 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2933__B key_in[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_402 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_785 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_424 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3748__C _3759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3110__A _3110_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_479 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_99 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_849 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5242__B1_N _5241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_859 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5037__A _4975_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_787 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_32 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4876__A _4876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3894__A2_N _3893_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3780__A _3780_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_223 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3106__A2 _3176_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_245 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4595__B _4595_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_671 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2865__A1 _2907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_343 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_900 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_977 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3202__A2_N _3201_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3020__A _3020_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5031__A2 _5017_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3955__A _5534_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_356 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4790__A1 _3231_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_602 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3847__A2_N _3846_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4790__B2 _4782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_304 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3674__B _3674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_808 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_540 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3393__C _5537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4370_ _4375_/A _4370_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_153_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_870 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_936 VGND VPWR sky130_fd_sc_hd__fill_1
X_3321_ _3320_/X _3321_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_724 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4786__A _3155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_81 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_958 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_3252_ _3110_/A _3251_/A _5497_/Q _3251_/Y _3253_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_86_619 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4845__A2 _4843_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_693 VGND VPWR sky130_fd_sc_hd__decap_12
X_3183_ _3116_/A _3183_/B _3185_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_121_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_719 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4058__B1 _4046_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_730 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4952__C _4951_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_251 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3281__A1 _3217_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5518__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_402 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_785 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_711 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4671__D _4670_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_424 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4026__A _4026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_435 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_109 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5022__A2 _5020_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1013 VGND VPWR sky130_fd_sc_hd__decap_6
X_2967_ _2966_/A _2965_/Y _2966_/X _2980_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3865__A _3861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_4706_ _2984_/A _4699_/X data_out2[14] _4701_/X _5416_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_120_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_507 VGND VPWR sky130_fd_sc_hd__decap_4
X_2898_ _2898_/A key_in[44] _2898_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_135_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3584__B _3584_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2792__B1 _2828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_635 VGND VPWR sky130_fd_sc_hd__decap_12
X_4637_ _4637_/A _4637_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3987__A1_N _3154_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_4568_ _4533_/X _4574_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_1_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_3519_ _3519_/A _2885_/A _5541_/Q _3519_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__4696__A _5522_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_532 VGND VPWR sky130_fd_sc_hd__fill_2
X_4499_ _4501_/A _4499_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_446 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5089__A2 _5087_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_479 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_332 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3105__A _5529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_343 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_985 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_996 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_23 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2944__A _2944_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_869 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5306__A2_N _5334_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3759__B _3758_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3272__B2 _3271_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_722 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_766 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_479 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_276 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3775__A _3773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_624 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_495 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_645 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3327__A2 _3324_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_3_0_clock_A clkbuf_4_3_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_188 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_595 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_405 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2838__B _2837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_62 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_84 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5486__RESET_B _4379_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3015__A _3015_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_803 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5415__RESET_B _4464_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_847 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2854__A _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_858 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_655 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5230__A _3608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_221 VGND VPWR sky130_fd_sc_hd__fill_2
X_3870_ _3870_/A _3869_/X _3870_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_32_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5004__A2 _4987_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_254 VGND VPWR sky130_fd_sc_hd__decap_3
X_2821_ _2741_/A _2799_/X _2752_/A _2799_/A _2799_/B _2821_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_32_788 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_290 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_991 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_440 VGND VPWR sky130_fd_sc_hd__fill_2
X_5540_ _3518_/X _5540_/Q _4314_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3566__A2 _2852_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_451 VGND VPWR sky130_fd_sc_hd__decap_12
X_2752_ _2752_/A _2801_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_76_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_635 VGND VPWR sky130_fd_sc_hd__decap_6
X_5471_ _5089_/X _5076_/A _4396_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_129_197 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_483 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_657 VGND VPWR sky130_fd_sc_hd__decap_12
X_4422_ _4422_/A _4422_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_711 VGND VPWR sky130_fd_sc_hd__fill_1
X_4353_ _4349_/A _4353_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_906 VGND VPWR sky130_fd_sc_hd__decap_8
X_3304_ _3304_/A _3304_/B _3304_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_59_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_928 VGND VPWR sky130_fd_sc_hd__fill_2
X_4284_ _4289_/A _4284_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_885 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2748__B _2745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_204 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5124__B _5114_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4666__D _4666_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_3235_ _3233_/X _3258_/A _3257_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_101_749 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2829__A1 _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_630 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_259 VGND VPWR sky130_fd_sc_hd__decap_12
X_3166_ _3143_/C _3166_/B _3166_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_493 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2764__A _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3097_ _3075_/Y _3095_/A _3096_/X _3099_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_54_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_655 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5140__A _5133_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_132 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_817 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3579__B _3577_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5497__D _5497_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_699 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_722 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_48 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_530 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5490__CLK _5430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_541 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_766 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_552 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_930 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_276 VGND VPWR sky130_fd_sc_hd__decap_8
X_3999_ _3939_/X _3998_/X _3999_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_22_287 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3595__A _3596_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_35 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_635 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4203__B _4203_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_808 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_370 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4857__C _4856_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4926__B1_N _4925_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_107 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5034__B _5031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_298 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4873__B _4872_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_825 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4690__B1 data_out2[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_644 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_99 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_869 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5050__A _5037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3489__B _3541_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_560 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_165 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_705 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3796__A2 _5527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_585 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_983 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4113__B _4113_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_475 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3952__B _3938_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2849__A _2849_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5225__A _5513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_928 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3720__A2 _3709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_939 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_758 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_180 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_257 VGND VPWR sky130_fd_sc_hd__fill_2
X_3020_ _3020_/A _3020_/B _3020_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_95_268 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_419 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_814 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_471 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4681__B1 data_out2[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_482 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_346 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3399__B _3398_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_4971_ _4971_/A _4970_/X _4971_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_64_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_338 VGND VPWR sky130_fd_sc_hd__fill_1
X_3922_ _3876_/Y _3922_/B _3922_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4984__A1 _5463_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_390 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_552 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2995__B1 _2958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_3853_ _3840_/Y _3852_/X _3853_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_2804_ _5198_/A _2772_/X _2736_/Y _2804_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4304__A _4304_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_900 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_207 VGND VPWR sky130_fd_sc_hd__decap_6
X_3784_ _3739_/Y _3783_/X _3759_/X _3785_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__2747__B1 _2746_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_781 VGND VPWR sky130_fd_sc_hd__decap_12
X_5523_ _5523_/D _5523_/Q _4335_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2735_ _2734_/Y _2735_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4023__B _4021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_123 VGND VPWR sky130_fd_sc_hd__decap_3
X_5454_ _4881_/X _4871_/A _4417_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4958__B _4958_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_318 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_273 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3862__B _3842_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4405_ _4419_/A _4411_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5161__A1 _5477_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_446 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2759__A _4882_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5385_ _4768_/X data_out1[15] _4499_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_530 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5135__A _5113_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4336_ _4339_/A _4336_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_563 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_725 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_224 VGND VPWR sky130_fd_sc_hd__decap_12
X_4267_ reset _4267_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4974__A _5463_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_3218_ _3145_/X key_in[53] _3218_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_825 VGND VPWR sky130_fd_sc_hd__decap_6
X_4198_ _4198_/A _4198_/B _4200_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_55_611 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3475__B2 _3474_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_3149_ _3145_/X key_in[115] _3044_/X _3149_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_43_806 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_463 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_23 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_725 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_596 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_747 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_900 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4727__A1 _3316_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4727__B2 _4726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4532__A1_N _4517_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2738__B1 _5287_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_944 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4868__B _4866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_424 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3772__B _3771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5386__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5152__A1 _5143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5045__A _5027_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4587__C _4578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_479 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3491__C _3490_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_874 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_682 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_622 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_482 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_817 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_891 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3012__B _3012_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_850 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_513 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2977__B1 _2937_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3947__B _3945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2851__B _2850_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_73 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_579 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_421 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3963__A _3958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_465 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3756__A1_N _2796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3154__B1 _3197_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_788 VGND VPWR sky130_fd_sc_hd__decap_6
X_5170_ _4891_/A _5170_/B _5170_/C _5170_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__5430__RESET_B _4445_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_170 VGND VPWR sky130_fd_sc_hd__fill_1
X_4121_ _4112_/X _4120_/Y _4123_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2901__B1 _2828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_490 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4794__A _3322_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_909 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_544 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_4052_ _3932_/Y _4048_/X _4051_/Y _4052_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_37_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_238 VGND VPWR sky130_fd_sc_hd__decap_6
X_3003_ _2968_/A key_in[111] _2828_/X _3003_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_110_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_806 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3203__A _3175_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_828 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_603 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_260 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4018__B _4018_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_327 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_113 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_967 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_809 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4957__B2 _4956_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4954_ _2973_/A _4954_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3709__A1_N _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3857__B _3812_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3905_ _3905_/A _3905_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_51_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_894 VGND VPWR sky130_fd_sc_hd__decap_4
X_4885_ _4885_/A _4884_/X _4885_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4709__A1 _5527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4709__B2 _4701_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3836_ data_in1[12] _3697_/X _3812_/X _3835_/Y _3836_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_165_538 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_3767_ _3701_/X _3709_/X _3766_/Y _3756_/X _3767_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_146_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_977 VGND VPWR sky130_fd_sc_hd__fill_2
X_5506_ _5506_/D _3251_/A _4355_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2718_ _2718_/A _2718_/B _2744_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_119_999 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5518__RESET_B _4341_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3698_ _4537_/X _3765_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_161_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_424 VGND VPWR sky130_fd_sc_hd__decap_3
X_5437_ _5437_/D _5203_/A _4437_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_10_69 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_254 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_608 VGND VPWR sky130_fd_sc_hd__fill_2
X_5368_ _2707_/A key_in[70] _5368_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_120_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_202 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3696__A1 data_in1[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4200__C _4200_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_298 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_833 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_170 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_4319_ _4340_/A _4324_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_5299_ _5299_/A _5300_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_59_268 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_599 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3448__B2 _3447_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_57 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_806 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3113__A _3113_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_901 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_934 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_33 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_411 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2952__A _2930_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5215__A1_N _5198_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4948__A1 _4943_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_308 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__B _3709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3620__A1 _3603_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_371 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3620__B2 _3603_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3555__A2_N _3554_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_527 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_538 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4879__A _4877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_599 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_432 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3783__A _3759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3384__B1 _3367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_231 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_788 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4884__B1 _4908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_674 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2846__B _2846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3439__B2 _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4119__A _4020_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_430 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_709 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3023__A _2997_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5401__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_293 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_669 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_455 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3072__C1 _3071_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_343 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5551__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4670_ _4527_/X _4616_/X _4661_/X _4669_/X _4670_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_159_387 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_229 VGND VPWR sky130_fd_sc_hd__fill_2
X_3621_ _5253_/Y _2734_/Y _3621_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_128_741 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3693__A _3694_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_508 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_774 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3914__A2 _3912_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3552_ _3529_/A key_in[95] _3552_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_722 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_744 VGND VPWR sky130_fd_sc_hd__fill_2
X_3483_ _3463_/Y _3482_/B _3540_/A _3489_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_131_906 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_608 VGND VPWR sky130_fd_sc_hd__fill_2
X_5222_ _5222_/A _5222_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_928 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4020__C _4019_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_118 VGND VPWR sky130_fd_sc_hd__decap_4
X_5153_ _5133_/Y _5147_/Y _5140_/B _5146_/X _5152_/X _5159_/A VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_97_864 VGND VPWR sky130_fd_sc_hd__fill_1
X_4104_ _4052_/X _4079_/X _4055_/Y _4104_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_111_663 VGND VPWR sky130_fd_sc_hd__fill_2
X_5084_ _5084_/A _5084_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_69_599 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2756__B key_in[72] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5132__B _5131_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4035_ _3848_/X _4011_/X _3999_/Y _4035_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4029__A _3905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_761 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_986 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3018__A1_N _2999_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_720 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4971__B _4970_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_113 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3850__B2 _3849_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_764 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3587__B _3587_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_797 VGND VPWR sky130_fd_sc_hd__decap_8
X_4937_ _4925_/X _4928_/X _4937_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3602__B2 _3590_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_842 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_825 VGND VPWR sky130_fd_sc_hd__decap_4
X_4868_ _4865_/X _4866_/X _4868_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_341 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_335 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4158__A2 _4154_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_730 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4699__A _4699_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3819_ _3819_/A _3797_/X _3819_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_165_357 VGND VPWR sky130_fd_sc_hd__fill_2
X_4799_ _5543_/Q _4799_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_20_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_774 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_936 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_593 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5307__B _5270_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5107__A1 _5104_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_232 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3108__A _3108_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3669__B2 _3668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_864 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4223__A2_N _3521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5323__A _5285_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5424__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4881__A3 _4880_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_374 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2892__A2 _2891_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_931 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_953 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_964 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_901 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_761 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5291__B1 _5325_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_986 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_485 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_76 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3841__A1 _3636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_945 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3841__B2 _3133_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5574__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_282 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3778__A _3778_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_753 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_455 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_978 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_168 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_691 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_831 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_663 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_149 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_97 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_875 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_886 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_869 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5346__B2 _5345_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_357 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_396 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4402__A _4402_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_1010 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5217__B _5216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4121__B _4120_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_906 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3109__B1 _3870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_928 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_980 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3960__B _3935_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2857__A _5358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_706 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_238 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_344 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4085__A1 _4784_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5282__B1 _5252_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_772 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_433 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_989 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_797 VGND VPWR sky130_fd_sc_hd__fill_2
X_2983_ _2998_/C _2982_/Y _2998_/C _2982_/Y _2984_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_691 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_296 VGND VPWR sky130_fd_sc_hd__decap_4
X_4722_ _5534_/Q _3287_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_195 VGND VPWR sky130_fd_sc_hd__decap_12
X_4653_ _4577_/A _4522_/A _4666_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_163_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_357 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3348__B1 _3333_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3604_ _5513_/Q _5518_/Q _3603_/X _3604_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__4312__A _4312_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_4584_ _4521_/A _4629_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_128_593 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4669__D _4668_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_221 VGND VPWR sky130_fd_sc_hd__decap_12
X_3535_ _3533_/X _3534_/Y _3533_/X _3534_/Y _3535_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4031__B _4030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_606 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5447__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_27 VGND VPWR sky130_fd_sc_hd__fill_1
X_3466_ _3155_/Y _3466_/B _3466_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_107_38 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4966__B _4965_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_49 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4946__A1_N _4553_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3260__B1_N _3305_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3870__B _3869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_758 VGND VPWR sky130_fd_sc_hd__decap_6
X_5205_ _4618_/A key_in[65] _5205_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2767__A _2767_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3397_ _5510_/Q _3397_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5143__A _5143_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_812 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_983 VGND VPWR sky130_fd_sc_hd__fill_1
X_5136_ _5110_/X _5137_/B _5136_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_85_823 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_37 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_5067_ _5566_/Q _5066_/X _5566_/Q _5066_/X _5067_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4982__A _4982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4076__A1 _3858_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4076__B2 _3463_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5273__B1 _5263_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_377 VGND VPWR sky130_fd_sc_hd__fill_1
X_4018_ _3966_/Y _4018_/B _4018_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_934 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_271 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_720 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_945 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3823__B2 _3822_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3110__B _3110_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5533__RESET_B _4323_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_847 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_67 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5318__A _5317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3339__B1 _3337_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_688 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_clock_A clkbuf_3_2_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_552 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_243 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_894 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4876__B _4874_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_736 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_66 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_521 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_235 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_514 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_471 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2865__A2 _2863_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_791 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_547 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2796__A1_N _2785_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_355 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5093__A1_N _5568_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4177__A2_N _4176_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_783 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_764 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5016__B1 _5562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_572 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_85 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3020__B _3020_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5031__A3 _5009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_611 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_632 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_171 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4790__A2 _4781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_120 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_143 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_154 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5228__A _5481_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_508 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_614 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_828 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_142 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__A _4000_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_316 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3971__A _3968_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3320_ _3320_/A _3320_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_153_883 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_224 VGND VPWR sky130_fd_sc_hd__decap_12
X_3251_ _3251_/A _3251_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_101_909 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_769 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_609 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4845__A3 _4844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3182_ _3160_/A _3182_/B _3182_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_66_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4058__B2 _4057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_366 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_837 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_347 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4307__A _4305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3211__A _3206_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3281__A2 _3280_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_926 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_948 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4026__B _3950_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_745 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5022__A3 _5021_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_2966_ _2966_/A _2965_/Y _2966_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3865__B _3864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4705_ _5525_/Q _2984_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_817 VGND VPWR sky130_fd_sc_hd__decap_3
X_2897_ _2896_/A _2895_/Y _2896_/X _2915_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_147_154 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5138__A _5138_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2792__A1 _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_102 VGND VPWR sky130_fd_sc_hd__decap_12
X_4636_ _4636_/A _4637_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_163_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_26 VGND VPWR sky130_fd_sc_hd__decap_4
X_4567_ _5568_/Q _4557_/B _4567_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_144_861 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_3518_ data_in2[29] _3391_/X _3493_/X _3517_/Y _3518_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_143_371 VGND VPWR sky130_fd_sc_hd__fill_1
X_4498_ _4501_/A _4498_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_393 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_544 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5089__A3 _5096_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_469 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_25 VGND VPWR sky130_fd_sc_hd__fill_2
X_3449_ _5473_/Q _3410_/X _3416_/X _3449_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_98_970 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_709 VGND VPWR sky130_fd_sc_hd__fill_1
X_5119_ _5129_/A _5118_/X _5129_/A _5118_/X _5119_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_355 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_804 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_34 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_163 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_clock_A clkbuf_3_5_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_314 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_325 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2944__B _2944_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_859 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_68 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4217__A _4215_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_959 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_266 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3152__B1_N _3196_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_644 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3775__B _3774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_809 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4887__A _4864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_541 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3167__B1_N _3166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_668 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3791__A _3780_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_894 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_853 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_81 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_7_0_clock_A clkbuf_4_7_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_812 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_823 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_739 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_791 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3015__B _2966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5237__B1 _5303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_51 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2854__B _2698_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_196 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5230__B _2716_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_358 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4127__A _4126_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5455__RESET_B _4416_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_241 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_166 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_211 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_408 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3966__A _3110_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2820_ _2819_/A _2819_/B _2872_/A _2822_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__2870__A _2870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_931 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_280 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_952 VGND VPWR sky130_fd_sc_hd__decap_12
X_2751_ _2750_/X _2752_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3566__A3 _5542_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_463 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_603 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_451 VGND VPWR sky130_fd_sc_hd__decap_6
X_5470_ _5075_/X _5470_/Q _4398_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_157_496 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4421_ _4422_/A _4421_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_466 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_861 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_872 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_894 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_371 VGND VPWR sky130_fd_sc_hd__fill_1
X_4352_ _4349_/A _4352_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_3303_ _3108_/Y _3303_/B _3304_/B VGND VPWR sky130_fd_sc_hd__nor2_4
X_4283_ _4304_/A _4289_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_255 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2748__C _5296_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3206__A _3135_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3234_ _3233_/A _3233_/B _3258_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_98_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2829__A2 key_in[106] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_642 VGND VPWR sky130_fd_sc_hd__decap_8
X_3165_ _3162_/X _3164_/Y _3162_/X _3164_/Y _3166_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_984 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_837 VGND VPWR sky130_fd_sc_hd__decap_6
X_3096_ _3073_/C _3096_/B _3096_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_81_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5140__B _5140_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_358 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_369 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3579__C _3596_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4037__A _4778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_520 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_205 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2780__A _2778_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_920 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_564 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3998_ _3903_/X _3964_/X _3952_/X _3987_/X _3998_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3595__B _3594_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2949_ _2998_/B _2948_/X _2998_/B _2948_/X _2989_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_806 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4203__C _4203_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4619_ _5236_/A _2707_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_2_605 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4500__A _4501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3201__A2_N _3200_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_406 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3116__A _3116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_750 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4690__A1 _5518_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5331__A _5331_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4690__B2 _4688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3846__A2_N _3845_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_336 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_756 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_391 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_542 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3786__A _3829_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_575 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_60 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_956 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_850 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4410__A _4411_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2849__B _2849_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_853 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3181__A1 _3180_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5508__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_341 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3026__A _3026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_374 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4130__B1 _3848_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_450 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4681__A1 _5513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5241__A _5239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_826 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_601 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_910 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4681__B2 _4677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_932 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_494 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2692__B1 _5356_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_976 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_464 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_550 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3986__A1_N _3984_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4970_ _4958_/X _4962_/X _4970_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_45_870 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_892 VGND VPWR sky130_fd_sc_hd__decap_4
X_3921_ _3873_/Y _3921_/B _3922_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_520 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4984__A2 _4847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2995__A1 data_in2[14] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_216 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_564 VGND VPWR sky130_fd_sc_hd__decap_12
X_3852_ _3875_/A _3850_/X _3851_/X _3852_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_20_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_238 VGND VPWR sky130_fd_sc_hd__fill_2
X_2803_ _2796_/X _2802_/X _2796_/X _2802_/X _2814_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_748 VGND VPWR sky130_fd_sc_hd__decap_8
X_3783_ _3759_/A _3758_/X _3783_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2747__A1 _5325_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5522_ _2882_/X _5522_/Q _4336_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3944__B1 _3943_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2734_ _2733_/C _2734_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_145_411 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_293 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_956 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_978 VGND VPWR sky130_fd_sc_hd__fill_2
X_5453_ _4869_/X _4859_/A _4418_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_157 VGND VPWR sky130_fd_sc_hd__decap_12
X_4404_ _4267_/Y _4419_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4320__A _4324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2759__B _2759_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5384_ _4766_/X data_out1[14] _4500_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5161__A2 _4995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_542 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5135__B _5135_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4335_ _4339_/A _4335_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_661 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3627__B1_N _3626_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_4266_ _4515_/A _4266_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_940 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_236 VGND VPWR sky130_fd_sc_hd__decap_12
X_3217_ _3217_/A _3212_/Y _3244_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5377__RESET_B _4508_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4197_ _4158_/X _4182_/B _4198_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_984 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_174 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_3148_ _3148_/A key_in[83] _3148_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_336 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_453 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4990__A _4978_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_3079_ _3043_/X key_in[113] _3044_/X _3079_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_54_166 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_998 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3632__C1 _3631_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_46 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_536 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_203 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4727__A2 _4725_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_923 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2738__A1 _5290_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2738__B2 _2943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_124 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_647 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_606 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_903 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_797 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_925 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4230__A _4794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_959 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5152__A2 _5145_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_831 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_458 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5045__B _5034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4587__D _4586_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_715 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_981 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_374 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4112__B1 _4786_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5061__A _5059_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_634 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_391 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_81 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2977__A1 _2905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_525 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3947__C _3947_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4405__A _4419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_884 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_96 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_591 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3963__B _3962_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_774 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5236__A _5236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3738__A2_N _3737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_105 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4140__A _4129_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3154__B2 _3153_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_650 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2901__A1 _2898_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4120_ _4114_/Y _4120_/B _4118_/Y _4119_/Y _4120_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_68_225 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5480__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_344 VGND VPWR sky130_fd_sc_hd__fill_2
X_4051_ _4050_/X _4051_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_110_366 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5470__RESET_B _4398_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_770 VGND VPWR sky130_fd_sc_hd__fill_2
X_3002_ _2790_/A key_in[79] _3002_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_37_634 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_667 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3203__B _3203_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_818 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_773 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_935 VGND VPWR sky130_fd_sc_hd__decap_8
X_4953_ _4943_/A _4847_/X _4942_/X _4952_/X _4953_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3614__C1 _3613_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_158 VGND VPWR sky130_fd_sc_hd__decap_6
X_3904_ _3794_/A _3903_/X _3904_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3857__C _3870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4315__A _4312_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4884_ _4908_/C _4883_/X _4908_/C _4883_/X _4884_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4709__A2 _4699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_534 VGND VPWR sky130_fd_sc_hd__decap_12
X_3835_ _3835_/A _3833_/Y _3834_/X _3835_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__2947__A2_N _2946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_422 VGND VPWR sky130_fd_sc_hd__decap_12
X_3766_ _3737_/X _3766_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_590 VGND VPWR sky130_fd_sc_hd__decap_12
X_5505_ _4166_/X _3231_/A _4356_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_146_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5244__A2_N _5243_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2717_ _2717_/A _2717_/B _2718_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_118_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_252 VGND VPWR sky130_fd_sc_hd__fill_2
X_3697_ _4533_/X _3697_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5146__A _5143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_488 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_274 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4050__A _4049_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_499 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_285 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_5436_ _4532_/X _5436_/Q _4438_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_127 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_458 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_469 VGND VPWR sky130_fd_sc_hd__decap_12
X_5367_ _2707_/A key_in[6] _5367_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4985__A _5464_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5558__RESET_B _4293_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4200__D _4200_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3696__A2 _3581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_523 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_823 VGND VPWR sky130_fd_sc_hd__fill_1
X_4318_ _4267_/Y _4340_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_5298_ _5234_/A _5299_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_19_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_355 VGND VPWR sky130_fd_sc_hd__decap_8
X_4249_ _4246_/X _4247_/Y _4248_/Y _4249_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_142_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_781 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_656 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3113__B _3088_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_637 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_45 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_423 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_283 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_125 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2952__B _2988_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4948__A2 _4946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_456 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_311 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4225__A _4225_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__C _3766_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_845 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_884 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3620__A2 _2723_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_681 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_709 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_366 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_377 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_505 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_388 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_55 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_591 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_77 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4879__B _4878_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3783__B _3758_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3384__B2 _3419_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_263 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5056__A _5056_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_200 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_734 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_722 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_766 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4895__A _5223_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3094__A2_N _3093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4884__B2 _4883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_276 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_545 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_409 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_515 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3304__A _3304_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_645 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4119__B _4119_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3023__B _3065_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_442 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_902 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_979 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3072__B1 _3026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_489 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3974__A _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3620_ _3603_/A _2723_/A _3619_/Y _3603_/X _3624_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3693__B _3692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4593__A1_N _5440_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_550 VGND VPWR sky130_fd_sc_hd__decap_3
X_3551_ _3529_/A key_in[31] _3551_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_701 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_3482_ _3463_/Y _3482_/B _3540_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_143_778 VGND VPWR sky130_fd_sc_hd__decap_8
X_5221_ _4529_/X _5222_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_5152_ _5143_/X _5145_/Y _5132_/Y _5152_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4103_ _4077_/X _4103_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_29_409 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_5083_ _5076_/Y _5079_/X _5082_/Y _5087_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_2_60 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3214__A _3170_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_239 VGND VPWR sky130_fd_sc_hd__decap_8
X_4034_ _3230_/X _4033_/X _3230_/X _4033_/X _4034_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_965 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4029__B _4028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_250 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_581 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_732 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5376__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_158 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3063__B1 _3074_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4045__A _4044_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4936_ _4642_/Y _4934_/X _4949_/A _4938_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
X_4867_ _4865_/X _4866_/X _4867_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_165_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3884__A _3823_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_325 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_859 VGND VPWR sky130_fd_sc_hd__fill_2
X_3818_ _2918_/A _3816_/X _3817_/X _3818_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_4798_ _5543_/Q _4798_/B _4798_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_2_3_0_clock_A clkbuf_2_3_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_561 VGND VPWR sky130_fd_sc_hd__decap_12
X_3749_ _3739_/Y _3744_/Y _3749_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_107_948 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5107__A2 _5103_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_918 VGND VPWR sky130_fd_sc_hd__decap_3
X_5419_ _5419_/D data_out2[17] _4459_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5392__RESET_B _4491_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_769 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5323__B _5322_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_984 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_729 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_921 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3124__A _3124_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_559 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5291__A1 _5290_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_913 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_464 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2963__A _2945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_529 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3841__A2 _5529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3778__B _3777_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_242 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_467 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_106 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_798 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_54 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_76 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3794__A _3794_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_825 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_364 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_38 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_807 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_745 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5409__RESET_B _4471_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3109__A1 _2961_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_541 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3109__B2 _3108_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_726 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_480 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3708__A1_N _3706_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2857__B _2887_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2868__B1 _5229_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_450 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_857 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5399__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_356 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5282__A1 data_in2[3] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4085__A2 _4083_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3969__A _3113_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_946 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_445 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_776 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2979__A1_N _2974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_938 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3045__B1 _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2982_ _2999_/A _2981_/X _2888_/Y _2982_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_15_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_681 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_139 VGND VPWR sky130_fd_sc_hd__fill_2
X_4721_ _4720_/X _4712_/X data_out2[22] _4713_/X _5424_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4793__B1 data_out1[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_314 VGND VPWR sky130_fd_sc_hd__fill_2
X_4652_ _4819_/A _4809_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_163_818 VGND VPWR sky130_fd_sc_hd__decap_3
X_3603_ _3603_/A _3603_/B _3603_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3348__B2 _3347_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_870 VGND VPWR sky130_fd_sc_hd__fill_1
X_4583_ _4582_/X _3465_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3209__A _3137_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3534_ _5143_/X _3504_/X _3507_/X _3534_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_155_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_564 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2917__A1_N _2888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_789 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_3465_ _3465_/A _3465_/B _3465_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_153_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_203 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5214__A1_N _5202_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_128 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_428 VGND VPWR sky130_fd_sc_hd__decap_8
X_5204_ _4618_/A key_in[1] _5204_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_640 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_247 VGND VPWR sky130_fd_sc_hd__fill_2
X_3396_ _3231_/Y _3396_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5135_ _5113_/A _5135_/B _5137_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_504 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_194 VGND VPWR sky130_fd_sc_hd__decap_12
X_5066_ _5037_/X _5065_/X _5066_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_879 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4982__B _4980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4076__A2 _5539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3879__A _3873_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_507 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5273__B2 _5272_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2783__A _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4017_ _4775_/X _3990_/X _4020_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_93_890 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_283 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_968 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_540 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_776 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_618 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_4919_ _4907_/A _4847_/X _4531_/X _4918_/X _4919_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_40_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_303 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4503__A _4501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3339__A1 _4639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_678 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_183 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5318__B _5317_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_194 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3339__B2 _3338_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_306 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_817 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_701 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_828 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5573__RESET_B _4274_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_892 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_839 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3119__A _3077_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_745 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5502__RESET_B _4359_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_361 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2958__A _3026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_715 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0_clock_A clkbuf_3_6_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5334__A _4836_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_383 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_940 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5541__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_312 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5264__A1 _4817_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_98 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_827 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_250 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_31 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_434 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_445 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5016__B2 _5015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_264 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_461 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_303 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4413__A _4418_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_110 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_154 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4132__B _4131_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3029__A _2999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3971__B _3970_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_916 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3017__A1_N _3892_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_61 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_512 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1000 VGND VPWR sky130_fd_sc_hd__decap_6
X_3250_ _4582_/X _3249_/X _3250_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_98_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_236 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_813 VGND VPWR sky130_fd_sc_hd__decap_4
X_3181_ _3180_/A _3180_/B _3236_/A _3187_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_94_610 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_559 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3699__A _3765_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_816 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_153 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_592 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_754 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_860 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3211__B _3210_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3018__B1 _2999_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_798 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4026__C _4778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_595 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_757 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_601 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4766__B1 data_out1[14] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2841__A1_N _2815_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2965_ _2944_/B _2965_/B _2964_/Y _2965_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_148_623 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_971 VGND VPWR sky130_fd_sc_hd__fill_1
X_4704_ _2989_/A _4699_/X data_out2[13] _4701_/X _5415_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4323__A _4324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5414__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2896_ _2896_/A _2895_/Y _2896_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_492 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_678 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5138__B _5138_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_4635_ _4635_/A _4636_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2792__A2 key_in[105] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_16 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_38 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5191__B1 _5182_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4566_ _4566_/A _4561_/B _4566_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_116_531 VGND VPWR sky130_fd_sc_hd__decap_12
X_3517_ _3317_/X _3517_/B _3517_/C _3517_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__2778__A _2778_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5564__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4497_ _4269_/A _4501_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5154__A _5477_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_748 VGND VPWR sky130_fd_sc_hd__fill_2
X_3448_ _5116_/A _3447_/X _5116_/A _3447_/X _3450_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_982 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4993__A _4985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_59 VGND VPWR sky130_fd_sc_hd__decap_3
X_3379_ _5472_/Q _3379_/B _3413_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_943 VGND VPWR sky130_fd_sc_hd__decap_3
X_5118_ _5037_/X _5129_/B _5118_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_643 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5246__A1 _3603_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_976 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_827 VGND VPWR sky130_fd_sc_hd__decap_4
X_5049_ _5469_/Q _5054_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_84_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3402__A _3400_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4217__B _4218_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_562 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_882 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_938 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_14_0_clock_A clkbuf_3_7_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3009__B1 _3050_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_921 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_960 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_623 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5329__A _5327_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4233__A _4230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_807 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_604 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_829 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5182__B1 _5181_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4887__B _4887_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3791__B _3786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_821 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5064__A _5470_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_692 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_865 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_556 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_919 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_898 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3496__B1 _3495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_470 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_654 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5237__A1 _5234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4408__A _4411_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_581 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2854__C _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3312__A _3312_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4127__B _4090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4003__B1_N _4002_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_882 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5437__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3966__B _3965_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2870__B _2870_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5495__RESET_B _4368_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_943 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VPWR sky130_fd_sc_hd__decap_3
X_2750_ _2742_/X _2749_/Y _2750_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_292 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3420__B1 _3320_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5424__RESET_B _4453_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_807 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_829 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_997 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3982__A _3858_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4420_ _4422_/A _4420_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_607 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_478 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_629 VGND VPWR sky130_fd_sc_hd__fill_1
X_4351_ _4349_/A _4351_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_692 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_320 VGND VPWR sky130_fd_sc_hd__fill_2
X_3302_ _3108_/Y _3303_/B _3304_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_4_691 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1019 VGND VPWR sky130_fd_sc_hd__fill_1
X_4282_ _4276_/X _4282_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_779 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_267 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3206__B _3209_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3233_ _3233_/A _3233_/B _3233_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_140_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_941 VGND VPWR sky130_fd_sc_hd__decap_12
X_3164_ _4582_/X _3163_/X _3107_/B _3164_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_67_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_518 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4318__A _4267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3239__B1 _3177_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3095_ _3095_/A _3096_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3222__A _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3524__A1_N _3396_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_808 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4037__B _4036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_702 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_871 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_882 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_908 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4739__B1 data_out2[31] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2780__B _2777_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3997_ _4026_/A _3950_/B _3010_/A _3997_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_22_256 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5149__A _5147_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_576 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4053__A _4002_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2948_ _4661_/X _2916_/Y _2888_/Y _2948_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3411__B1 _5473_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_604 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_818 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4988__A _4985_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2879_ _2855_/Y _2921_/B _2879_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_129_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3892__A _3892_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4176__A2_N _4175_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4618_ _4618_/A _5236_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_840 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_884 VGND VPWR sky130_fd_sc_hd__decap_12
X_4549_ _5552_/Q _4541_/B _4549_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_132_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_556 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3116__B _3115_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_898 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_654 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_451 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_762 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4690__A2 _4687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_540 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_819 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_189 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3786__B _3785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5059__A _5059_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_72 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_935 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_412 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_434 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5155__B1 _5144_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_455 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_372 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3181__A2 _3180_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_353 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3026__B _2884_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4130__A1 _4096_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_676 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_985 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4681__A2 _4674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5241__B _5241_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_922 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_838 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4138__A _4788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_944 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2692__B2 _2691_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3042__A _2861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_540 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_988 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3977__A _4537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2881__A _2852_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3920_ _3872_/Y _3896_/Y _3920_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4884__A1_N _4908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_690 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2995__A2 _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3851_ _3875_/A _3850_/X _3851_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_2802_ _2802_/A _2801_/X _2802_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_81_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_751 VGND VPWR sky130_fd_sc_hd__decap_12
X_3782_ _3743_/X _3782_/B _3831_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_5521_ _2853_/X _5521_/Q _4337_/X _5402_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3944__A1 _2889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2747__A2 _5332_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2733_ _2733_/A _2698_/B _2733_/C _2733_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_157_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_794 VGND VPWR sky130_fd_sc_hd__decap_6
X_5452_ _5452_/D _4848_/A _4420_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4601__A _5443_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_242 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_478 VGND VPWR sky130_fd_sc_hd__fill_2
X_4403_ _4402_/A _4403_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_169 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_938 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_489 VGND VPWR sky130_fd_sc_hd__fill_2
X_5383_ _4764_/X data_out1[13] _4501_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3217__A _3217_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_843 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_459 VGND VPWR sky130_fd_sc_hd__decap_4
X_4334_ _4339_/A _4334_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_716 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_898 VGND VPWR sky130_fd_sc_hd__decap_6
X_4265_ _4629_/D _4264_/B all_done _5434_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_86_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_3216_ _3216_/A _3143_/B _4718_/X _3216_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4196_ _4156_/X _4196_/B _4196_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_28_816 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_304 VGND VPWR sky130_fd_sc_hd__fill_1
X_3147_ _3077_/A key_in[19] _3147_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_82_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_635 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_819 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_605 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4990__B _4983_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3078_ _3077_/A key_in[81] _3078_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_860 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_638 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2791__A _2898_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3632__B1 _3615_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_852 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_863 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_716 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_885 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_548 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_896 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2738__A2 _2737_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_434 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_220 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_136 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4511__A _4269_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_916 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4230__B _4212_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_425 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3127__A _3048_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_959 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_843 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_180 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_993 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_161 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2966__A _2966_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_56 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5342__A _4848_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4112__B2 _4111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5061__B _5058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_985 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_827 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3797__A _3682_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_627 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_649 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3623__B1 _5272_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_532 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2977__A2 _2976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_42 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_537 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_902 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_743 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4421__A _4422_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_905 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_776 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5236__B key_in[66] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4140__B _4159_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_437 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3037__A _3014_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_662 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_215 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2901__A2 key_in[108] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2876__A _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5252__A _5252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_194 VGND VPWR sky130_fd_sc_hd__decap_12
X_4050_ _4049_/X _4050_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_451 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_218 VGND VPWR sky130_fd_sc_hd__fill_2
X_3001_ _2790_/A key_in[15] _3001_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_49_473 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5402__D _5402_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_495 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4193__A1_N _4187_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_955 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_741 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_657 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_292 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_977 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_465 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_4952_ _4918_/A _4950_/X _4951_/Y _4952_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3614__B1 _3599_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3500__A _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3903_ _3884_/X _3893_/X _3903_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4883_ _4874_/A _4872_/X _4873_/A _4883_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_32_384 VGND VPWR sky130_fd_sc_hd__decap_12
X_3834_ _3827_/X _3832_/Y _3834_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_546 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_209 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_913 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3917__A1 _3904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_3765_ _3765_/A _3679_/B _3778_/A _3765_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_158_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_434 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4331__A _4330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5119__B1 _5129_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5504_ _4143_/X _3178_/A _4357_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2716_ _2716_/A _2717_/B _2718_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_3696_ data_in1[6] _3581_/X _3679_/X _3695_/X _3696_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_161_702 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_404 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5146__B _5145_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_798 VGND VPWR sky130_fd_sc_hd__decap_3
X_5435_ _5435_/D _4256_/A _4439_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_10_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_5366_ _5299_/A key_in[38] _5366_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_373 VGND VPWR sky130_fd_sc_hd__fill_2
X_4317_ _4312_/A _4317_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2786__A _5300_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5297_ _5294_/A _5294_/B _5325_/B _5297_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_59_237 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_868 VGND VPWR sky130_fd_sc_hd__decap_6
X_4248_ _5197_/A _3788_/A _5510_/Q data_in1[31] _4546_/A _4248_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_142_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_613 VGND VPWR sky130_fd_sc_hd__fill_2
X_4179_ _4791_/X _4177_/X _4196_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_55_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_281 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5527__RESET_B _4330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_668 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3605__B1 _5242_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4506__A _4504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_830 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_301 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_874 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4225__B _4224_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__D _3756_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_334 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_693 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_879 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_170 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_34 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_517 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_34 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_89 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5337__A _2707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_701 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_651 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4895__B _4918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_778 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2696__A _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_288 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_621 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_632 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3688__B1_N _3687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5072__A _5072_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_194 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_602 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3304__B _3304_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_527 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_624 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_955 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4416__A _4418_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3320__A _3320_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_159 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3072__A1 data_in2[16] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_991 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3308__A1_N _3290_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5349__B1 _5321_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_367 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_866 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_209 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3974__B _3972_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_754 VGND VPWR sky130_fd_sc_hd__decap_4
X_3550_ _3528_/A key_in[63] _3550_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_127_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_562 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_275 VGND VPWR sky130_fd_sc_hd__decap_12
X_3481_ _3465_/Y _3480_/Y _3465_/Y _3480_/Y _3482_/B VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_170_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_757 VGND VPWR sky130_fd_sc_hd__fill_2
X_5220_ data_in2[1] _4574_/B _5197_/X _5219_/X _5220_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_115_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_256 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2897__B1_N _2896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_418 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_470 VGND VPWR sky130_fd_sc_hd__decap_12
X_5151_ _4857_/A _5149_/X _5150_/Y _5143_/X _4815_/A _5476_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_97_855 VGND VPWR sky130_fd_sc_hd__fill_2
X_4102_ _3980_/Y _4098_/X _4101_/Y _4102_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_111_654 VGND VPWR sky130_fd_sc_hd__fill_2
X_5082_ _5081_/X _5082_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_911 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2820__B1_N _2872_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_387 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3214__B _3212_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4033_ _4031_/X _4032_/X _4031_/X _4032_/X _4033_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_72 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_432 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_752 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_413 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4326__A _4340_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_744 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3063__A1 _3062_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_660 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4045__B _4034_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4935_ _4642_/Y _4934_/X _4949_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_833 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_310 VGND VPWR sky130_fd_sc_hd__fill_2
X_4866_ _4852_/X _4855_/X _4866_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_21_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3154__A2_N _3153_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3884__B _3847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_877 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_710 VGND VPWR sky130_fd_sc_hd__fill_1
X_3817_ _2918_/A _3816_/X _3817_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4797_ _5510_/Q _4674_/A data_out1[31] _4677_/A _4797_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4012__B1 _3999_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5147__B1_N _5146_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4061__A _4072_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3748_ _3765_/A _3679_/B _3759_/A _3748_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_137_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_787 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4996__A _4996_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3679_ _3615_/A _3679_/B _4750_/X _3679_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_118_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_19 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_459 VGND VPWR sky130_fd_sc_hd__decap_8
X_5418_ _4709_/X data_out2[16] _4460_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_256 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_971 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_610 VGND VPWR sky130_fd_sc_hd__fill_2
X_5349_ _5321_/C _5348_/X _5321_/C _5348_/X _5351_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_470 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_332 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3405__A _3337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_654 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_974 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_741 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5291__A2 _5290_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_605 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2963__B _2944_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_700 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_733 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4236__A _3676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3140__A _3139_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3737__A2_N _3736_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_11 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_254 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_788 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_84 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_811 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_118 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_991 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_310 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_321 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_676 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_332 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_804 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5470__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_88 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_815 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3794__B _3793_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_175 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_849 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_376 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_819 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_540 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_871 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_882 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_554 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3109__A2 _3108_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_418 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_597 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2868__A1 _2717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2868__B2 _3032_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5449__RESET_B _4423_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3315__A _5355_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_85 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_335 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_741 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5282__A2 _5222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_903 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3969__B _3942_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2946__A2_N _2945_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5243__A2_N _5242_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_593 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4146__A _3394_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_232 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3050__A _2974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_906 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_917 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3045__A1 _3043_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2981_ _2998_/A _2998_/B _2981_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4242__B1 _4731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4793__A1 _3300_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4720_ _4720_/A _4720_/X VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4793__B2 _4677_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_849 VGND VPWR sky130_fd_sc_hd__decap_12
X_4651_ _4651_/A _4819_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_3602_ _3588_/Y _3589_/Y _3573_/X _3590_/X _3619_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4582_ _2999_/A _4582_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3209__B _3209_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3533_ _5154_/Y _3532_/Y _5154_/Y _3532_/Y _3533_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_746 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_3464_ _3464_/A _3464_/B _3465_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_103_418 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_373 VGND VPWR sky130_fd_sc_hd__fill_2
X_5203_ _5203_/A key_in[33] _5203_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_930 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_321 VGND VPWR sky130_fd_sc_hd__fill_2
X_3395_ _3394_/Y _3395_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_630 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3225__A _5468_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_652 VGND VPWR sky130_fd_sc_hd__decap_8
X_5134_ _5134_/A _5122_/A _5138_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_29_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_387 VGND VPWR sky130_fd_sc_hd__decap_8
X_5065_ _5065_/A _5051_/X _5065_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4016_ _3968_/X _4019_/B _4016_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3879__B _3877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2783__B _2698_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_947 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_733 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4056__A _4052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_232 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5493__CLK _5430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_939 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_585 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3895__A _3895_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_4918_ _4918_/A _4916_/Y _4917_/X _4918_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_139_827 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_315 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_47 VGND VPWR sky130_fd_sc_hd__decap_12
X_4849_ _5547_/Q _4838_/B _4849_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_138_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_696 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3339__A2 _3335_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_860 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3119__B key_in[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2958__B _2884_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_727 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5334__B _5334_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_790 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3135__A _3069_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_952 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5542__RESET_B _4312_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_836 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5350__A _5350_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_806 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5264__A2 _5238_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_763 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_305 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_402 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_593 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5500__D _4042_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4224__B1 _4207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_438 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_473 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_674 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3029__B _3028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_690 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_521 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_862 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_939 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_524 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_215 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_790 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_3180_ _3180_/A _3180_/B _3236_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_836 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_538 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2884__A _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_110 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5260__A _5260_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_132 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_806 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_666 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3699__B _3679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_165 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5410__D _5410_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_552 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_574 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3018__B2 _3017_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_980 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4766__A1 _3870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4766__B2 _4758_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2964_ _2896_/A _2964_/B _2895_/Y _2964_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_4703_ _5524_/Q _2989_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_123 VGND VPWR sky130_fd_sc_hd__decap_4
X_2895_ _2871_/B _2893_/Y _2894_/Y _2895_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_136_808 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_60 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_605 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5138__C _5136_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4634_ _4616_/X _4633_/X _2907_/A _4616_/X _5437_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_871 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_126 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3442__B1_N _3441_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4565_ _5566_/Q _4561_/B _5566_/D VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__5191__B2 _5190_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_874 VGND VPWR sky130_fd_sc_hd__fill_2
X_3516_ _3516_/A _3516_/B _3517_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2778__B _2777_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4496_ _4492_/A _4496_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_513 VGND VPWR sky130_fd_sc_hd__decap_12
X_3447_ _4640_/X _3443_/X _3444_/X _3445_/X _3446_/X _3447_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_131_579 VGND VPWR sky130_fd_sc_hd__decap_8
X_3378_ _4639_/X _3374_/X _3375_/X _3376_/X _3377_/X _3379_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_57_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_922 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_782 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2794__A _5456_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_5117_ _5569_/Q _5101_/X _5129_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_281 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5170__A _4891_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5246__A2 _5245_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5048_ _4896_/X _5046_/Y _5047_/X _5036_/Y _4806_/X _5048_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_84_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_560 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3402__B _3401_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1011 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_917 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_799 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4206__B1 _4073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3009__B2 _3008_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_900 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4514__A _4515_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_35 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2768__B1 _2767_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_972 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5329__B _5327_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_635 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4233__B _4233_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_616 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_189 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5389__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5182__A1 _3578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2969__A _2934_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5345__A _2769_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_863 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3193__B1 _3191_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_800 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_65 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3496__A1 _4788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_611 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4693__B1 data_out2[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_397 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5080__A _5076_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5237__A2 key_in[98] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_64 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3312__B _3352_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_658 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_755 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_97 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4127__C _4788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_703 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_179 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4424__A _4422_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_8 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_972 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_271 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_955 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_282 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3420__A1 _3465_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_293 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_189 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3982__B _3981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_435 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2879__A _2855_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5255__A _5227_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5464__RESET_B _4406_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4350_ _4349_/A _4350_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_362 VGND VPWR sky130_fd_sc_hd__decap_4
X_3301_ _3158_/A _3300_/A _4775_/X _3466_/B _3303_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_4281_ _4276_/X _4281_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5405__D _4682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_888 VGND VPWR sky130_fd_sc_hd__decap_12
X_3232_ _2889_/Y _3231_/A _3113_/A _3231_/Y _3233_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_39_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_398 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_482 VGND VPWR sky130_fd_sc_hd__fill_2
X_3163_ _3028_/X _3163_/B _3163_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_95_953 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_997 VGND VPWR sky130_fd_sc_hd__fill_2
X_3094_ _3176_/B _3093_/X _3176_/B _3093_/X _3095_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3239__A1 _4661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_474 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_647 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_360 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4739__A1 _5542_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4334__A _4339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4739__B2 _4737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_911 VGND VPWR sky130_fd_sc_hd__decap_4
X_3996_ data_in1[19] _3976_/X _3978_/X _3995_/Y _5498_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_22_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5149__B _5149_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_27 VGND VPWR sky130_fd_sc_hd__fill_2
X_2947_ _2939_/X _2946_/X _2939_/X _2946_/X _2998_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4053__B _4029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3411__B2 _3410_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5531__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_791 VGND VPWR sky130_fd_sc_hd__fill_2
X_2878_ _2878_/A _2920_/B _2921_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4988__B _4987_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_947 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3892__B _3891_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4617_ _5203_/A _4618_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2789__A _2790_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_969 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_468 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5165__A _5165_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_351 VGND VPWR sky130_fd_sc_hd__decap_4
X_4548_ _4908_/C _4547_/B _4548_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_896 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_4479_ _4477_/A _4479_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_257 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4124__C1 _4123_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_568 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3478__A1 _3475_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4509__A _4504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_953 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3413__A _3340_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_552 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3016__A1_N _3036_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_533 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3646__A1_N _3635_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4244__A _4244_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_257 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5059__B _5058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_599 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_55 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1003 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_785 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_402 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_947 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_638 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_649 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5155__A1 _4572_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_969 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_446 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2699__A _2885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_979 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_811 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_833 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_408 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3026__C _5527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_899 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_611 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_920 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_92 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4130__A2 _4109_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_249 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4419__A _4419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3917__B1_N _3916_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5404__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4851__A2_N _4850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_997 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4138__B _4137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_625 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3042__B key_in[80] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4969__A1 _3052_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_563 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2881__B _2879_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_371 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5554__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_382 VGND VPWR sky130_fd_sc_hd__fill_2
X_3850_ _3847_/X _3849_/X _3847_/X _3849_/X _3850_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_886 VGND VPWR sky130_fd_sc_hd__decap_3
X_2801_ _2801_/A _2801_/B _2801_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_739 VGND VPWR sky130_fd_sc_hd__decap_3
X_3781_ _3778_/A _3777_/X _3828_/A _3829_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_13_791 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3993__A _3979_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_240 VGND VPWR sky130_fd_sc_hd__decap_4
X_5520_ _2811_/X _5520_/Q _4338_/X _5402_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_118_605 VGND VPWR sky130_fd_sc_hd__decap_4
X_2732_ _5223_/A _2733_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_30_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3944__A2 _3941_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_402 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_273 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_947 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_272 VGND VPWR sky130_fd_sc_hd__decap_3
X_5451_ _4845_/X _4836_/A _4421_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4601__B _4601_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_906 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_928 VGND VPWR sky130_fd_sc_hd__decap_4
X_4402_ _4402_/A _4402_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_800 VGND VPWR sky130_fd_sc_hd__decap_12
X_5382_ _5382_/D data_out1[12] _4502_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_427 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_833 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3217__B _3212_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4333_ _4340_/A _4339_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_577 VGND VPWR sky130_fd_sc_hd__decap_4
X_4264_ _4662_/Y _4264_/B _4264_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_101_505 VGND VPWR sky130_fd_sc_hd__decap_12
X_3215_ data_in2[20] _3172_/X _3174_/X _3214_/Y _5531_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4329__A _4330_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4195_ _3466_/B _4193_/Y _4231_/A _4195_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_79_290 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_132 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3233__A _3233_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_901 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_603 VGND VPWR sky130_fd_sc_hd__decap_6
X_3146_ _3145_/X key_in[51] _3146_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_95_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_124 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_967 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_3077_ _3077_/A key_in[17] _3077_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_872 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_488 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3632__A1 data_in1[3] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4064__A _4778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_363 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_739 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_227 VGND VPWR sky130_fd_sc_hd__decap_6
X_3979_ _3966_/Y _3972_/Y _3979_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5386__RESET_B _4498_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_468 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3408__A _3222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_416 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3127__B _3127_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_437 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_855 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_674 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5427__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2966__B _2965_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5342__B _5341_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_441 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3143__A _3026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_997 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_400 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4647__B1_N _4646_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_95 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5577__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_669 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5073__B1 _4803_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3797__B _3796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4820__B1 _4541_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3623__B2 _3622_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_10 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_330 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_886 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_897 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_914 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_273 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_703 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3318__A _3318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_736 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_991 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_286 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3037__B _3037_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_503 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2876__B _2876_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_696 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_324 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5252__B _5252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3538__A1_N _3521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_869 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4149__A _4147_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3000_ _2898_/A key_in[47] _3000_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_49_463 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_783 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_422 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3988__A _3903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1003 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_230 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_499 VGND VPWR sky130_fd_sc_hd__decap_8
X_4951_ _4951_/A _4949_/X _4951_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_17_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_959 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3614__A1 data_in1[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_842 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3500__B key_in[61] VGND VPWR sky130_fd_sc_hd__diode_2
X_3902_ _3839_/A _3812_/B _3902_/C _3902_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4882_ _4882_/A _4885_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_503 VGND VPWR sky130_fd_sc_hd__decap_12
X_3833_ _3827_/X _3832_/Y _3833_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_20_525 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3378__B1 _3376_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_903 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_558 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3917__A2 _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_925 VGND VPWR sky130_fd_sc_hd__fill_2
X_3764_ data_in1[9] _3697_/X _3748_/X _3763_/Y _5488_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_158_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_5503_ _5503_/D _3155_/A _4358_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5119__B2 _5118_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2715_ _3626_/A _2714_/A _5260_/A _2714_/Y _2717_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_446 VGND VPWR sky130_fd_sc_hd__decap_6
X_3695_ _3676_/A _3693_/X _3694_/Y _3695_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3228__A _5023_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5434_ _5434_/D all_done _4441_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_133_416 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_5365_ _5364_/A _5363_/Y _5364_/X _5365_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_160_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_983 VGND VPWR sky130_fd_sc_hd__decap_12
X_4316_ _4312_/A _4316_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5362__B1_N _2719_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_825 VGND VPWR sky130_fd_sc_hd__decap_8
X_5296_ _5296_/A _5325_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4059__A _4043_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4247_ _4246_/A _4246_/B _3579_/A _4247_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_68_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_923 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3384__A2_N _3419_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_4178_ _4791_/X _4177_/X _4178_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_68_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_891 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_647 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3898__A _3883_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_3129_ _3129_/A _3127_/X _3128_/Y _3129_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_76_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_14 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5055__B1 _5072_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_477 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_628 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_105 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3605__B2 _3604_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_436 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_803 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5567__RESET_B _4282_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_661 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_503 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_672 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_374 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_346 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_508 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_547 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3369__B1 _4778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_46 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4522__A _4522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5337__B key_in[5] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5315__B1_N _5350_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_435 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3138__A _3135_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_713 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_980 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4869__B1 _4859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5353__A _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_994 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2696__B _2694_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5072__B _5072_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_569 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5503__D _5503_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_60 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3601__A _3586_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_488 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_959 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3072__A2 _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_801 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_335 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5349__B2 _5348_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_160 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_182 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3974__C _3973_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_711 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4432__A _4426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_878 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_221 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3048__A _3048_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3480_ _3469_/X _3479_/X _3469_/X _3479_/X _3480_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_142_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_544 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2887__A _2887_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3532__B1 _3530_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5150_ _5147_/Y _5149_/B _5150_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_111_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_482 VGND VPWR sky130_fd_sc_hd__decap_6
X_4101_ _4100_/X _4101_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_5081_ _5080_/X _5081_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_867 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_121 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5413__D _5413_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_677 VGND VPWR sky130_fd_sc_hd__decap_4
X_4032_ _4002_/X _4009_/X _4032_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_99_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_260 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3214__C _3213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_444 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4607__A _4609_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_455 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_978 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3511__A _3493_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_105 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_937 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_425 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_778 VGND VPWR sky130_fd_sc_hd__decap_4
X_4934_ _4944_/A _4933_/X _4944_/A _4933_/X _4934_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3063__A2 _3061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4045__C _3998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_683 VGND VPWR sky130_fd_sc_hd__fill_2
X_4865_ _4863_/A _4862_/X _4864_/Y _4865_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_60_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_867 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4342__A _4341_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3816_ _2735_/X _5528_/Q _2733_/C _3075_/Y _3816_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_20_344 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3884__C _3866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_891 VGND VPWR sky130_fd_sc_hd__fill_2
X_4796_ _3368_/A _4674_/A data_out1[30] _4677_/A _4796_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4012__B2 _4011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_3747_ data_in1[8] _3697_/X _3719_/X _3746_/Y _3747_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_21_38 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_928 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3771__B1 _5356_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_939 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_416 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_3678_ _4664_/X _3679_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_134_747 VGND VPWR sky130_fd_sc_hd__fill_1
X_5417_ _4708_/X data_out2[15] _4461_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2797__A _2797_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_268 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5173__A _5355_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5348_ _5324_/Y _5347_/Y _5324_/Y _5347_/Y _5348_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_153_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_738 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3405__B key_in[26] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_5279_ _5277_/X _5280_/B _5281_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_75_506 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_753 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4517__A _5436_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_639 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4236__B _4236_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3140__B _3138_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_767 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_650 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_622 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_288 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_171 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_480 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_806 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_817 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_688 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_519 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_344 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4252__A _4576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_699 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4003__A1 _3175_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_349 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_850 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_232 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_359 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_500 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4192__A1_N _3479_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_265 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_823 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_460 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_739 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_920 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_42 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2868__A2 _3902_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_953 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_355 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_804 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_506 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_97 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_377 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_314 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5489__RESET_B _4375_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4427__A _4426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5418__RESET_B _4460_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3331__A _3331_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_745 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4146__B _4145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3050__B _3050_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3045__A2 key_in[112] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4242__A1 _4047_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2980_ _2980_/A _2980_/B _2998_/C VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__4242__B2 _3548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_672 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_620 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4793__A2 _4674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5258__A _5258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_165 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4162__A _4159_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4650_ _4524_/A _4650_/B _4518_/A _4649_/X _4651_/A VGND VPWR sky130_fd_sc_hd__or4_4
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_338 VGND VPWR sky130_fd_sc_hd__decap_12
X_3601_ _3586_/A _3600_/X _3601_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__5408__D _4689_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4581_ _5358_/A _2999_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_360 VGND VPWR sky130_fd_sc_hd__fill_2
X_3532_ _4640_/X _3528_/X _3529_/X _3530_/X _3531_/X _3532_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_155_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_909 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_769 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_706 VGND VPWR sky130_fd_sc_hd__fill_2
X_3463_ _5539_/Q _3463_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_408 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3505__B1 _5143_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5202_ _5181_/X _5201_/X _5181_/X _5201_/X _5202_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_739 VGND VPWR sky130_fd_sc_hd__fill_2
X_3394_ _5537_/Q _3394_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_130_238 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3225__B _3226_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5133_ _5132_/A _5131_/X _5132_/Y _5133_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_96_130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_986 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_697 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_5064_ _5470_/Q _5068_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_731 VGND VPWR sky130_fd_sc_hd__decap_12
X_4015_ _3972_/A _4015_/B _4019_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_37_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4337__A _4339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_369 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_775 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2783__C _2847_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3241__A _4718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_937 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_414 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3672__B1_N _3671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4056__B _4055_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_907 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_981 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3895__B _3894_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_597 VGND VPWR sky130_fd_sc_hd__decap_3
X_4917_ _4917_/A _4915_/Y _4917_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_15 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5168__A _5169_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2795__A1 _4900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_625 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_839 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4072__A _4072_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4848_ _4848_/A _4852_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_21_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_59 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_48 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3339__A3 _3336_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4779_ _4778_/X _4769_/X data_out1[21] _4770_/X _4779_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_153_319 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4800__A _4799_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4941__C1 _4940_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_831 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3610__B1_N _3595_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_596 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_544 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_886 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2958__C _2984_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3416__A _3416_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3135__B _3099_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_964 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3307__A1_N _3299_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_152 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_196 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5350__B _5319_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_230 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_904 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_509 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_818 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3151__A _5013_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5511__RESET_B _4349_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_892 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_745 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_66 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4224__A1 _4000_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_981 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4224__B2 _4209_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_597 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_299 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5078__A _5037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_951 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_485 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_973 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_658 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_668 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_168 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4710__A _5528_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_544 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_841 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3326__A _3325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_85 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_569 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_848 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_794 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2884__B _2884_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_196 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4157__A _4156_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3699__C _5229_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_572 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_417 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_439 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4766__A2 _4757_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2963_ _2945_/A _2944_/A _2965_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_31_940 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2777__A1 _2723_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4702_ _5523_/Q _4699_/X data_out2[12] _4701_/X _5414_/D VGND VPWR sky130_fd_sc_hd__o22a_4
X_2894_ _2822_/A _2871_/X _2821_/X _2894_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_129_850 VGND VPWR sky130_fd_sc_hd__decap_4
X_4633_ _3529_/A _4631_/Y _4800_/B _4631_/A _4633_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__5138__D _5137_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_72 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3726__B1 _3725_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4620__A _2707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_680 VGND VPWR sky130_fd_sc_hd__decap_12
X_4564_ _5065_/A _4561_/B _4564_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_149 VGND VPWR sky130_fd_sc_hd__decap_4
X_3515_ _3516_/A _3516_/B _3517_/B VGND VPWR sky130_fd_sc_hd__nor2_4
X_4495_ _4492_/A _4495_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_171_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3236__A _3236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_525 VGND VPWR sky130_fd_sc_hd__fill_1
X_3446_ _3499_/A key_in[123] _3408_/X _3446_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_131_536 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4151__B1 _3417_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3377_ _3334_/X key_in[121] _3222_/X _3377_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_58_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_472 VGND VPWR sky130_fd_sc_hd__fill_2
X_5116_ _5116_/A _5121_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_85_623 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5460__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2794__B _2794_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_336 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_956 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5170__B _5170_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4067__A _4068_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_509 VGND VPWR sky130_fd_sc_hd__fill_1
X_5047_ _5047_/A _5045_/X _5047_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_27_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4206__A1 _4187_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_372 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_247 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2768__A1 _5334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3965__B1 _3954_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_450 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_422 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_984 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4233__C _4232_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_967 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_605 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4530__A _4529_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5182__A2 _3671_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2969__B key_in[14] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_649 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_853 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3193__A1 _4638_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5345__B _5345_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3193__B2 _3192_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_19 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3146__A _3145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_897 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_599 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_940 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2985__A _2984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_409 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4693__A1 _2847_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3496__A2 _4794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_77 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5361__A _5361_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4693__B2 _4688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_794 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5080__B _5079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5511__D _5196_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_54 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3653__C1 _3652_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_840 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_862 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4705__A _5525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_361 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_288 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_236 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_250 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__B1 _2984_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_411 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_283 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_995 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3420__A2 _3419_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_967 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_294 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_483 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_977 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3708__B1 _3706_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4440__A _4419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_447 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2879__B _2921_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5255__B _5254_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3056__A _2911_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_374 VGND VPWR sky130_fd_sc_hd__fill_2
X_3300_ _3300_/A _3466_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_514 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5483__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_396 VGND VPWR sky130_fd_sc_hd__fill_2
X_4280_ _4276_/X _4280_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_247 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_3231_ _3231_/A _3231_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2895__A _2871_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3092__A2_N _3091_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_377 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5433__RESET_B _4442_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_111 VGND VPWR sky130_fd_sc_hd__decap_12
X_3162_ _3154_/X _3161_/X _3154_/X _3161_/X _3162_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_591 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_965 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5421__D _5421_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3093_ _4582_/X _3060_/A _3060_/X _3093_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3239__A2 _3201_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4615__A _4629_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_726 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4739__A2 _4736_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3995_ _3974_/A _3993_/Y _3994_/X _3995_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_22_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_409 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_945 VGND VPWR sky130_fd_sc_hd__fill_2
X_2946_ _2964_/B _2945_/X _2964_/B _2945_/X _2946_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_967 VGND VPWR sky130_fd_sc_hd__fill_1
X_2877_ _2876_/A _2876_/B _2920_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_30_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_403 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4350__A _4349_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4616_ _4615_/X _4616_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_680 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2789__B key_in[9] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5165__B _5164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4547_ _4874_/A _4547_/B _5550_/D VGND VPWR sky130_fd_sc_hd__or2_4
Xclkbuf_4_13_0_clock clkbuf_3_6_0_clock/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_150_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_514 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_385 VGND VPWR sky130_fd_sc_hd__fill_1
X_4478_ _4477_/A _4478_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4124__B1 _4091_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3429_ _3426_/X _3429_/B _3431_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3478__A2 _3477_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5181__A _3577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_965 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3413__B _3413_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4525__A _4524_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_383 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_692 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_236 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4244__B _4243_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_567 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_720 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_910 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_230 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1015 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5356__A _5252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4260__A _4616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5155__A2 _5052_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5506__D _5506_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_300 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_653 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5091__A _4566_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_932 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4969__A2 _4968_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4435__A _4438_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_361 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2881__C _2880_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_821 VGND VPWR sky130_fd_sc_hd__decap_3
X_2800_ _2799_/A _2799_/B _2799_/X _2802_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
X_3780_ _3780_/A _3828_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3993__B _4015_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_2731_ _5222_/A _2731_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_904 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_797 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5266__A _5236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_211 VGND VPWR sky130_fd_sc_hd__decap_6
X_5450_ _4835_/X _4827_/A _4422_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_157_285 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4170__A _4152_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_447 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4401_ _4402_/A _4401_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_406 VGND VPWR sky130_fd_sc_hd__fill_2
X_5381_ _4761_/X data_out1[11] _4503_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5416__D _5416_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_812 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_439 VGND VPWR sky130_fd_sc_hd__decap_4
X_4332_ _4330_/A _4332_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1011 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_631 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_567 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_867 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_878 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_4263_ _4261_/X _4263_/B _4258_/C _4263_/D _4263_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_86_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_517 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3514__A _3540_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_932 VGND VPWR sky130_fd_sc_hd__decap_8
X_3214_ _3170_/A _3212_/Y _3213_/X _3214_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_4194_ _3466_/B _4193_/Y _4231_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3233__B _3233_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3145_ _3043_/X _3145_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_67_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_840 VGND VPWR sky130_fd_sc_hd__fill_1
X_3076_ _3043_/X key_in[49] _3076_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5379__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4345__A _4341_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3093__B1 _3060_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_681 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3632__A2 _3581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_534 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4064__B _4036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_38 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_353 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_729 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4042__C1 _4041_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3978_ _4026_/A _3950_/B _4775_/X _3978_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_50_375 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4593__B1 _5440_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_701 VGND VPWR sky130_fd_sc_hd__fill_1
X_2929_ _2733_/A _2884_/B _2989_/A _2929_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5176__A _5355_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_756 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_609 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_789 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_266 VGND VPWR sky130_fd_sc_hd__decap_12
X_5579_ _4264_/X _4518_/A _4266_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_491 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_366 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_377 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_68 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3424__A _3484_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_954 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3856__C1 _3855_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_41 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3143__B _3143_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5073__A1 _5071_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_979 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4255__A _4631_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3084__B1 _3128_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_990 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4820__B2 _4819_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_394 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_876 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_66 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_77 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_550 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_926 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_751 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_414 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_458 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3318__B _3318_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_748 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_683 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3505__A2_N _3504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3037__C _3036_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_826 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3334__A _3291_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_983 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5252__C _5514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4149__B _4149_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5521__CLK _5402_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_626 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3380__B1_N _3413_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3988__B _3964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1015 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_445 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4139__B1_N _4138_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4165__A _4092_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4950_ _4951_/A _4949_/X _4950_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_17_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_798 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_681 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_117 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3614__A2 _3581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_383 VGND VPWR sky130_fd_sc_hd__decap_12
X_3901_ data_in1[15] _3837_/X _3882_/X _3900_/Y _5494_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_32_320 VGND VPWR sky130_fd_sc_hd__decap_12
X_4881_ _4870_/X _4879_/Y _4880_/X _4871_/A _4815_/X _4881_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_60_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_353 VGND VPWR sky130_fd_sc_hd__decap_12
X_3832_ _3804_/X _3832_/B _3830_/Y _3831_/Y _3832_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_20_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_898 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3378__A1 _4639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3378__B2 _3377_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_561 VGND VPWR sky130_fd_sc_hd__fill_2
X_3763_ _3788_/A _3761_/Y _3762_/X _3763_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_5502_ _4089_/X _3108_/A _4359_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2714_ _2714_/A _2714_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_69_1005 VGND VPWR sky130_fd_sc_hd__decap_12
X_3694_ _3694_/A _3692_/X _3694_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3228__B _3228_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_778 VGND VPWR sky130_fd_sc_hd__decap_12
X_5433_ _4739_/X data_out2[31] _4442_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_156_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_5364_ _5364_/A _5363_/Y _5364_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_353 VGND VPWR sky130_fd_sc_hd__decap_12
X_4315_ _4312_/A _4315_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_815 VGND VPWR sky130_fd_sc_hd__decap_8
X_5295_ _5294_/X _5296_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_142_995 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3645__A1_N _5311_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3244__A _3244_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_325 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_16 VGND VPWR sky130_fd_sc_hd__fill_2
X_4246_ _4246_/A _4246_/B _4246_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__5026__A2_N _5025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4059__B _4058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_913 VGND VPWR sky130_fd_sc_hd__decap_3
X_4177_ _4171_/Y _4176_/Y _4171_/Y _4176_/Y _4177_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_870 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3898__B _3921_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3128_ _3128_/A _3128_/B _3057_/Y _3128_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_83_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5055__A1 _5054_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_905 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_916 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_253 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4075__A _4073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_489 VGND VPWR sky130_fd_sc_hd__fill_2
X_3059_ _3039_/X _3058_/X _3039_/X _3058_/X _3060_/B VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_36_670 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_949 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_297 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_448 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_815 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_459 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_640 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_353 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_898 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4803__A _4656_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_397 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3369__A1 _3233_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3369__B2 _3368_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_14 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_583 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3419__A _3419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5536__RESET_B _4320_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_745 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3138__B _3137_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_575 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4869__A1 _4802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_737 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4869__B2 _4815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_246 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5353__B _5351_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_130 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5544__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2696__C _2695_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_792 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_483 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2993__A _3065_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_946 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_99 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_968 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_220 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3601__B _3600_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4254__C1 _4253_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2804__B1 _2736_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_314 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_662 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_971 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_813 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4713__A _4701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_364 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_347 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_172 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3329__A _3259_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_380 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_531 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_778 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_789 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_748 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_556 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2887__B _2887_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5119__A1_N _5129_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3532__A1 _4640_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3532__B2 _3531_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3064__A _3064_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_537 VGND VPWR sky130_fd_sc_hd__decap_12
X_4100_ _4099_/X _4100_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_5080_ _5076_/Y _5079_/X _5080_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_133 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_667 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3999__A _3939_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4031_ _4029_/X _4030_/Y _4031_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_65_710 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_916 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3511__B _3539_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_949 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_437 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4796__B1 data_out1[30] VGND VPWR sky130_fd_sc_hd__diode_2
X_4933_ _4921_/X _4932_/X _4933_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_33_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_459 VGND VPWR sky130_fd_sc_hd__decap_6
X_4864_ _4863_/X _4864_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_60_470 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4623__A _2861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5417__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_334 VGND VPWR sky130_fd_sc_hd__fill_2
X_3815_ _3794_/A _3814_/X _3815_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_165_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3884__D _3814_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_356 VGND VPWR sky130_fd_sc_hd__decap_12
X_4795_ _4794_/X _4674_/A data_out1[29] _4677_/A _5399_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_165_339 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_391 VGND VPWR sky130_fd_sc_hd__decap_6
X_3746_ _3788_/A _3744_/Y _3745_/X _3746_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_118_233 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3771__A1 _3589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_501 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3771__B2 _3770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_715 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5567__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3677_ data_in1[5] _3581_/X _3654_/X _3676_/X _3677_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_118_288 VGND VPWR sky130_fd_sc_hd__decap_6
X_5416_ _5416_/D data_out2[14] _4463_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_115_951 VGND VPWR sky130_fd_sc_hd__decap_12
X_5347_ _5333_/X _5346_/X _5333_/X _5346_/X _5347_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_130_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_601 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_835 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_27 VGND VPWR sky130_fd_sc_hd__fill_2
X_5278_ _5278_/A _5278_/B _5280_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_87_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_667 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_518 VGND VPWR sky130_fd_sc_hd__fill_2
X_4229_ _3523_/X _4228_/X _3523_/X _4228_/X _4229_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3702__A _3681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_957 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_968 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_478 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_404 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_724 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_584 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4236__C _4236_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_297 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4787__B1 data_out1[24] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_64 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_267 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_982 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4533__A _4529_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_835 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_166 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_356 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3537__A1_N _3522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4003__A2 _4001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_839 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5370__RESET_B _4516_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2988__A _2925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_512 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5364__A _5364_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_567 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_718 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4711__B1 data_out2[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_577 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5514__D _5514_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_323 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_943 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_879 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_442 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_965 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_816 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3278__B1 _3354_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__A _3609_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_348 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3331__B _3330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_916 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4112__A2_N _4111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_949 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_256 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4242__A2 _5542_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5458__RESET_B _4413_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_982 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4443__A _4443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_306 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4162__B _4198_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_3600_ _3600_/A _3592_/Y _3600_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_128_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_4580_ _5256_/A _5358_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3202__B1 _3177_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3383__A2_N _3382_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_873 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3753__A1 _3636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3531_ _3528_/A key_in[126] _3408_/X _3531_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__2898__A _2898_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_883 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5274__A _5274_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_3462_ _3519_/A _3364_/B _5539_/Q _3462_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_5201_ _5199_/Y _5361_/A _3583_/C _5200_/A _5201_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4702__B1 data_out2[12] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3505__B2 _3504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_3393_ _3519_/A _3364_/B _5537_/Q _3393_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5424__D _5424_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_5132_ _5132_/A _5131_/X _5132_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_69_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_453 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_827 VGND VPWR sky130_fd_sc_hd__decap_12
X_5063_ _5469_/Q _4995_/X _4942_/X _5062_/X _5063_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4618__A _4618_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_4014_ _3180_/A _4012_/X _4013_/Y _4014_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_38_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_562 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3241__B _3280_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_724 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_437 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_565 VGND VPWR sky130_fd_sc_hd__fill_2
X_4916_ _4917_/A _4915_/Y _4916_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__4353__A _4349_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_481 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2795__A2 _2794_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3992__A1 _4775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5168__B _5169_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_654 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4072__B _4069_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4847_ _4891_/A _4847_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_4778_ _3030_/A _4778_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_361 VGND VPWR sky130_fd_sc_hd__decap_8
X_3729_ _3728_/X _3730_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_4_308 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4941__B1 _4531_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4800__B _4800_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_737 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5184__A _4618_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3416__B _3415_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4820__A1_N _4541_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_589 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3135__C _3068_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_131 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_431 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_751 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_475 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4528__A _4614_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3432__A _3317_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_551 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3151__B _3195_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_212 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_554 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4224__A2 _4097_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5359__A _5490_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_89 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5551__RESET_B _4301_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_587 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4263__A _4261_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_941 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5078__B _5077_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_637 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5509__D _5509_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_512 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5094__A _5090_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_853 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_567 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_504 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_352 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_886 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_762 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_613 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4438__A _4438_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2884__C _5523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3117__B1_N _3116_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_348 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_294 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4999__B1 _4559_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_562 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_584 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_830 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_297 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_757 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_971 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_716 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4173__A _4146_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2962_ _2961_/A _2961_/B _3015_/A _2966_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_97_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2777__A2 _2723_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4701_ _4701_/A _4701_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_963 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5419__D _5419_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_974 VGND VPWR sky130_fd_sc_hd__fill_2
X_2893_ _2872_/A _2871_/A _2893_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_147_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_4632_ _4798_/B _4800_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_129_862 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3726__A1 _2735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_84 VGND VPWR sky130_fd_sc_hd__decap_8
X_4563_ _5564_/Q _4557_/B _4563_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_129_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_692 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_680 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3517__A _3317_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3514_ _3540_/A _3491_/B _3516_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_545 VGND VPWR sky130_fd_sc_hd__decap_12
X_4494_ _4492_/A _4494_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3236__B _3187_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_3445_ _3501_/A key_in[91] _3445_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4634__A2_N _4633_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_559 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4151__B2 _4150_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_3376_ _3337_/A key_in[89] _3376_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_58_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_602 VGND VPWR sky130_fd_sc_hd__decap_8
X_5115_ _5473_/Q _4995_/X _4942_/X _5114_/Y _5115_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_58_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_175 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4348__A _4349_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_635 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5170__C _5170_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_5046_ _5047_/A _5045_/X _5046_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_73_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_27 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4067__B _4066_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_768 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4206__A2 _4192_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_15 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5179__A _3577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_15 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2768__A2 _2769_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3965__B2 _3964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_648 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_462 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4811__A _4811_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_350 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3427__A _4728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3193__A2 _3189_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3146__B key_in[51] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_762 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4693__A2 _4687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_366 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_827 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5361__B _5361_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4258__A _4252_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_370 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3653__B1 _3633_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_50 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_373 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_941 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_240 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__A1 _3750_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_963 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_259 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_262 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__B2 _3955_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_273 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_423 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_284 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_411 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_295 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_979 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_793 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_70 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_489 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3708__B2 _3707_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3337__A _3337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_342 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_705 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_650 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_727 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3056__B _3055_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_749 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_537 VGND VPWR sky130_fd_sc_hd__decap_12
X_3230_ _3227_/X _3229_/X _3227_/X _3229_/X _3230_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4133__A1 _4000_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_879 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2895__B _2893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_900 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4168__A _4157_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3161_ _3183_/B _3160_/X _3183_/B _3160_/X _3161_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_977 VGND VPWR sky130_fd_sc_hd__decap_4
X_3092_ _3937_/A _3091_/X _3937_/A _3091_/X _3176_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5473__RESET_B _4394_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_115 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3644__B1 _3666_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_830 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3800__A _3799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_841 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5402__RESET_B _4479_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4615__B _4615_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_738 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_3994_ _3979_/Y _4015_/B _3994_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_167_209 VGND VPWR sky130_fd_sc_hd__fill_2
X_2945_ _2945_/A _2896_/X _2945_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_148_434 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3306__A1_N _3304_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4631__A _4631_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2876_ _2876_/A _2876_/B _2878_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_148_478 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_415 VGND VPWR sky130_fd_sc_hd__decap_12
X_4615_ _4629_/B _4615_/B _4615_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3247__A _3216_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4546_ _4546_/A _4547_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3580__C1 _3579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_364 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_993 VGND VPWR sky130_fd_sc_hd__decap_12
X_4477_ _4477_/A _4477_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_237 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4124__A1 data_in1[24] VGND VPWR sky130_fd_sc_hd__diode_2
X_3428_ _3366_/A _3427_/X _3385_/X _3429_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_131_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5181__B _5181_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4078__A _3955_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3359_ _3359_/A _3359_/B _3357_/Y _3358_/Y _3359_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_85_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_732 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_454 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_860 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_988 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_871 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_5029_ _5027_/A _5027_/B _5028_/Y _5034_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4806__A _4815_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_532 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3710__A _3702_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_922 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4541__A _4541_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_765 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_927 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5356__B _2698_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_926 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_117 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4260__B _4659_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3157__A _3158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_469 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_982 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_898 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2996__A _3026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_481 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_492 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4083__A1_N _4075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5312__B1 _5297_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_507 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_664 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5091__B _5077_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5522__D _2882_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_830 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_874 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_524 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_833 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_170 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_192 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_731 VGND VPWR sky130_fd_sc_hd__fill_1
X_2730_ data_in2[7] _5222_/X _2698_/X _2729_/Y _5518_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4451__A _4449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5450__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4036__A1_N _4034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_415 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5266__B key_in[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_106 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4170__B _4136_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3067__A _2988_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_285 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_128 VGND VPWR sky130_fd_sc_hd__fill_2
X_4400_ _4402_/A _4400_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_60_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_5380_ _4759_/X data_out1[10] _4505_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_154_982 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_109 VGND VPWR sky130_fd_sc_hd__decap_12
X_4331_ _4330_/A _4331_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_992 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_491 VGND VPWR sky130_fd_sc_hd__decap_4
X_4262_ _4631_/Y _4654_/Y _4263_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_708 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_3213_ _3213_/A _3211_/X _3213_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3514__B _3491_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3314__C1 _3313_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_186 VGND VPWR sky130_fd_sc_hd__decap_12
X_4193_ _4187_/Y _4192_/Y _4187_/Y _4192_/Y _4193_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_68_944 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5432__D _5432_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_966 VGND VPWR sky130_fd_sc_hd__decap_12
X_3144_ _3144_/A _3139_/Y _3169_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_95_763 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_988 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_498 VGND VPWR sky130_fd_sc_hd__fill_2
X_3075_ _5528_/Q _3075_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4626__A _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3230__A1_N _3227_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_649 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3530__A _3529_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3093__A1 _4582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_340 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_660 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_991 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_181 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_490 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_507 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_708 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4042__B1 _4026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_888 VGND VPWR sky130_fd_sc_hd__fill_2
X_3977_ _4537_/X _4026_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_387 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4361__A _4267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_2928_ data_in2[12] _2731_/X _2884_/X _2927_/Y _5523_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_149_765 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4593__B2 _4590_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_253 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_927 VGND VPWR sky130_fd_sc_hd__fill_2
X_2859_ _2859_/A key_in[43] _2859_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_156_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_919 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_907 VGND VPWR sky130_fd_sc_hd__decap_4
X_5578_ _4263_/X _4522_/A _4271_/A _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_813 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_470 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_610 VGND VPWR sky130_fd_sc_hd__fill_1
X_4529_ _4528_/X _4529_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3705__A _2723_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5192__A _5178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5395__RESET_B _4487_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_849 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3856__B1 _3839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_421 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_890 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3143__C _3143_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_273 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4536__A _4529_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_424 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3440__A _3399_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5073__A2 _5072_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4255__B _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3084__B2 _3083_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_896 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_170 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_34 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5473__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4033__B1 _4031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5367__A _2707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3091__A2_N _3090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_61 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4271__A _4271_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_562 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5517__D _5517_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_734 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_982 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_952 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3615__A _3615_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_229 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2725__B1_N _2694_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_590 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3847__B1 _2939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_498 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_649 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4446__A _4443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_254 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_777 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4165__B _4168_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_822 VGND VPWR sky130_fd_sc_hd__decap_4
X_3900_ _3835_/A _3898_/Y _3899_/X _3900_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_17_395 VGND VPWR sky130_fd_sc_hd__decap_12
X_4880_ _4877_/X _4878_/X _4880_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5349__A1_N _5321_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_3831_ _3831_/A _3829_/X _3831_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_32_365 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3059__A2_N _3058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3378__A2 _3374_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4181__A _4168_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_398 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3689__A2_N _3688_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3762_ _3749_/Y _3782_/B _3762_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_158_551 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_550 VGND VPWR sky130_fd_sc_hd__fill_2
X_5501_ _4070_/X _3085_/A _4360_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2713_ _2704_/X _2712_/X _2704_/X _2712_/X _2713_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3693_ _3694_/A _3692_/X _3693_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5427__D _5427_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_768 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_705 VGND VPWR sky130_fd_sc_hd__decap_3
X_5432_ _5432_/D data_out2[30] _4443_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_215 VGND VPWR sky130_fd_sc_hd__decap_8
X_5363_ _5325_/X _5332_/A _5331_/A _5363_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_160_248 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_4314_ _4312_/A _4314_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5294_ _5294_/A _5294_/B _5294_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_462 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3244__B _3244_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4245_ _4239_/X _4244_/X _4239_/X _4244_/X _4246_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_229 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_538 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_730 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_605 VGND VPWR sky130_fd_sc_hd__decap_6
X_4176_ _3452_/X _4175_/X _3452_/X _4175_/X _4176_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_67_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_700 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_413 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_733 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_593 VGND VPWR sky130_fd_sc_hd__fill_2
X_3127_ _3048_/A _3127_/B _3127_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4356__A _4354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_295 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5055__A2 _5054_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5496__CLK _5429_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_766 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_928 VGND VPWR sky130_fd_sc_hd__decap_4
X_3058_ _3128_/A _3057_/Y _3128_/A _3057_/Y _3058_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4075__B _4074_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_118 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_827 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_315 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_849 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_365 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_337 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4091__A _4026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3369__A2 _3368_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_702 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_415 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3419__B _3419_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_971 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_418 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4869__A2 _4867_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_726 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5576__RESET_B _4271_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_749 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_790 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3435__A _3435_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5353__C _5352_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5505__RESET_B _4356_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_903 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2993__B _2991_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_893 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_649 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4266__A _4515_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_40 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_381 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3170__A _3170_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_906 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_608 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4254__B1 _4809_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_170 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2804__A1 _5198_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_674 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_899 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_825 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__A _5098_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_359 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_871 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3329__B _3304_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_212 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_746 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_520 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_768 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_593 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_705 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_92 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_597 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3345__A _3268_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_568 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3532__A2 _3528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3064__B _3020_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_357 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_291 VGND VPWR sky130_fd_sc_hd__fill_2
X_4030_ _3905_/Y _4028_/X _4030_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5273__A1_N _5263_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3999__B _3998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_722 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_969 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4245__B1 _4239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_671 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_276 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4910__A2_N _4909_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4904__A _4914_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4932_ _5554_/Q _4922_/X _4932_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4796__A1 _3368_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4796__B2 _4677_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4863_ _4863_/A _4862_/X _4863_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_847 VGND VPWR sky130_fd_sc_hd__decap_6
X_3814_ _3793_/X _3802_/X _3814_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4794_ _3322_/A _4794_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_702 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_368 VGND VPWR sky130_fd_sc_hd__decap_12
X_3745_ _3740_/X _3742_/X _3745_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_9_391 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3771__A2 _3020_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3676_ _3676_/A _3674_/X _3675_/Y _3676_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_118_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_5415_ _5415_/D data_out2[13] _4464_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_115_963 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_140 VGND VPWR sky130_fd_sc_hd__fill_2
X_5346_ _5335_/X _5345_/X _5335_/X _5345_/X _5346_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_707 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_985 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_922 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_112 VGND VPWR sky130_fd_sc_hd__fill_2
X_5277_ _5253_/Y _5276_/B _5276_/X _5277_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_101_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_988 VGND VPWR sky130_fd_sc_hd__decap_12
X_4228_ _4222_/X _4227_/X _4222_/X _4227_/X _4228_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_925 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_402 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_593 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3702__B _3701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4086__A _4072_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4159_ _4112_/X _4159_/B _4120_/Y _4159_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_83_541 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_619 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_788 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3039__A1 _3038_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_596 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4787__A1 _4786_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4814__A _4813_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4787__B2 _4782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_257 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_803 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2798__B1 _5327_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_814 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_302 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_306 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3747__C1 _3746_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_543 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5511__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_705 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2988__B _2988_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_512 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5364__B _5363_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3691__A1_N _4750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4711__A1 _3073_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4711__B2 _4701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_589 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_977 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3278__A1 _4720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__B _3610_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_733 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5530__D _3171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_530 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2713__A2_N _2712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_703 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_563 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4227__B1 _3535_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_630 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4724__A _5535_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_994 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_808 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_791 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_318 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_666 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5498__RESET_B _4365_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3202__B2 _3201_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_91 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5427__RESET_B _4450_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3753__A2 _3751_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3530_ _3529_/A key_in[94] _3530_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2898__B key_in[44] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__A1_N _3588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_895 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_738 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5274__B _5274_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_372 VGND VPWR sky130_fd_sc_hd__fill_2
X_3461_ data_in2[27] _3391_/X _3434_/X _3460_/Y _5538_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_171_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3075__A _5528_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_5200_ _5200_/A _5361_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4702__A1 _5523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4702__B2 _4701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_600 VGND VPWR sky130_fd_sc_hd__fill_2
X_3392_ _5223_/A _3519_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_922 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2713__B1 _2704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_622 VGND VPWR sky130_fd_sc_hd__decap_8
X_5131_ _5571_/Q _5130_/X _5571_/Q _5130_/X _5131_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_421 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5290__A _5290_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_508 VGND VPWR sky130_fd_sc_hd__decap_12
X_5062_ _4918_/A _5060_/Y _5061_/X _5062_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_96_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_839 VGND VPWR sky130_fd_sc_hd__decap_12
X_4013_ _3180_/A _4012_/X _4013_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_37_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5440__D _4593_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_287 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_298 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_449 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_769 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_577 VGND VPWR sky130_fd_sc_hd__decap_3
X_4915_ _4900_/X _4913_/X _4914_/X _4915_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_21_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_791 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5534__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_819 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3992__A2 _3990_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4846_ _4803_/Y _4891_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_165_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_841 VGND VPWR sky130_fd_sc_hd__decap_12
X_4777_ _3010_/A _4769_/X data_out1[20] _4770_/X _4777_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_119_532 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_705 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4941__A1 _4642_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3728_ _3728_/A _3685_/X _3706_/X _3728_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_10_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_885 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_502 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_576 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_896 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5184__B key_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_215 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_321 VGND VPWR sky130_fd_sc_hd__fill_2
X_3659_ _3588_/Y _5521_/Q _3588_/Y _5521_/Q _3659_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_899 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3901__C1 _3900_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_5329_ _5327_/A _5327_/B _5330_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4809__A _4799_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_443 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_817 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_677 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_999 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4528__B _4527_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_880 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_176 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_487 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3432__B _3432_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5103__A1_N _5569_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_872 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_13 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4209__B1 _4188_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_522 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4544__A _5548_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_769 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_57 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_268 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_419 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4263__B _4263_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_471 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_622 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_633 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_121 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_666 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2999__A _2999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_114 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_699 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_852 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5520__RESET_B _4338_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_351 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5094__B _5093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_693 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_855 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5525__D _5525_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_365 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_622 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_549 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_281 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_292 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5407__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_519 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_828 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_530 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4999__B2 _4998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_254 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5557__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4957__A1_N _4554_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4454__A _4449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_728 VGND VPWR sky130_fd_sc_hd__decap_4
X_2961_ _2961_/A _2961_/B _3015_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4173__B _4173_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_482 VGND VPWR sky130_fd_sc_hd__fill_2
X_4700_ _4700_/A _4701_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_1019 VGND VPWR sky130_fd_sc_hd__fill_1
X_2892_ _2714_/Y _2891_/B _2945_/A _2896_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_31_986 VGND VPWR sky130_fd_sc_hd__decap_12
X_4631_ _4631_/A _4631_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5285__A _5256_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_496 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3726__A2 _3722_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2702__A _5357_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4562_ _5563_/Q _4557_/B _4562_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3517__B _3517_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3513_ _3513_/A _3516_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_7_692 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_332 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5435__D _5435_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4493_ _4492_/A _4493_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_408 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_140 VGND VPWR sky130_fd_sc_hd__decap_12
X_3444_ _3501_/A key_in[27] _3444_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_171_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_3375_ _3337_/A key_in[25] _3375_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4629__A _4518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_817 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_903 VGND VPWR sky130_fd_sc_hd__fill_2
X_5114_ _4891_/A _5114_/B _5114_/C _5114_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_69_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_947 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3536__A1_N _3527_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_647 VGND VPWR sky130_fd_sc_hd__decap_12
X_5045_ _5027_/X _5034_/X _5045_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_27_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_703 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_725 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_680 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4364__A _4367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_875 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_925 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_49 VGND VPWR sky130_fd_sc_hd__fill_2
X_4829_ _4542_/A _4828_/X _4542_/A _4828_/X _4830_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_474 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4811__B _4810_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5195__A _5281_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_833 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3427__B _3385_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3193__A3 _3190_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_866 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_825 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4678__B1 data_out2[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_430 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4539__A _5197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_741 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_879 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3443__A _3499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_452 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_975 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3350__B1 _3320_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_603 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_251 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_262 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4258__B _4615_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_530 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_541 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_157 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_606 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3382__A2_N _3381_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_511 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3653__A1 data_in1[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_747 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_758 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4274__A _4271_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_886 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3956__A2 _5534_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_263 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_947 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_60 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_159 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3618__A _3586_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_416 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_822 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3337__B key_in[88] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_739 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_695 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4133__A2 _4131_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__A _4449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_194 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3965__A2_N _3964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2895__C _2894_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3353__A _3353_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_912 VGND VPWR sky130_fd_sc_hd__decap_3
X_3160_ _3160_/A _3116_/X _3160_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4168__B _4168_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_102 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_658 VGND VPWR sky130_fd_sc_hd__fill_2
X_3091_ _3112_/B _3090_/X _3112_/B _3090_/X _3091_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_308 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3644__A1 _3641_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_371 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_680 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_650 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_706 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_875 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_514 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_3993_ _3979_/Y _4015_/B _3993_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_149_903 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5442__RESET_B _4431_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2944_ _2944_/A _2944_/B _2964_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_936 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_906 VGND VPWR sky130_fd_sc_hd__decap_12
X_2875_ _2857_/Y _2887_/B _2857_/Y _2887_/B _2876_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_19 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3528__A _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4614_ _4525_/X _4629_/D _4614_/C _4615_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_135_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3247__B _3143_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_844 VGND VPWR sky130_fd_sc_hd__decap_6
X_4545_ _4545_/A _4541_/B _4545_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_117_855 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3580__B1 _3570_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_825 VGND VPWR sky130_fd_sc_hd__fill_2
X_4476_ _4469_/A _4477_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_132_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4359__A _4354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4124__A2 _3976_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3427_ _4728_/X _3385_/B _3427_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_89_249 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3263__A _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_912 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3475__A1_N _5128_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3358_ _3210_/Y _3357_/B _3358_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_38_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_411 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4078__B _4076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_593 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_669 VGND VPWR sky130_fd_sc_hd__decap_8
X_3289_ _3249_/X _3273_/X _3318_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_5028_ _5027_/X _5028_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_72_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_894 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_511 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3710__B _3709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_544 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4094__A _4073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_525 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_711 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_413 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_260 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4541__B _4541_/B VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_clock clkbuf_4_7_0_clock/A _5402_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3438__A _3465_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5356__C _5356_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_989 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4260__C _4255_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3157__B _3158_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_471 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2996__B _2884_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_633 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5312__B2 _5311_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4269__A _4269_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3173__A _5223_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3323__B1 _3010_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_208 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_923 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_422 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_179 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_469 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_801 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_783 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_794 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_293 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4170__C _4093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3067__B _3066_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_909 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_297 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_960 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3274__A2_N _3273_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4330_ _4330_/A _4330_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_674 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_493 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4179__A _4791_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4261_ _4629_/B _4522_/A _4615_/B _4261_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_113_346 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3314__B1 _3287_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3212_ _3213_/A _3211_/X _3212_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_113_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_4192_ _3479_/X _4191_/X _3479_/X _4191_/X _4192_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_95_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_433 VGND VPWR sky130_fd_sc_hd__fill_2
X_3143_ _3026_/A _3143_/B _3143_/C _3143_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_67_444 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4907__A _4907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_978 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5067__B1 _5566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3811__A _4664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_786 VGND VPWR sky130_fd_sc_hd__decap_3
X_3074_ _3074_/A _3071_/B _3099_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_54_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_680 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3530__B key_in[94] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3093__A2 _3060_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_867 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4642__A _4642_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3976_ _4533_/X _3976_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4042__A1 data_in1[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_2927_ _2927_/A _2925_/Y _2926_/X _2927_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3258__A _3258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_265 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_17 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_736 VGND VPWR sky130_fd_sc_hd__decap_12
X_2858_ _2858_/A _2838_/X _2858_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_145_950 VGND VPWR sky130_fd_sc_hd__fill_2
X_5577_ _4260_/X _4521_/A _4270_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2789_ _2790_/A key_in[9] _2789_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3553__B1 _3408_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4528_ _4614_/C _4527_/X _4528_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_117_685 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_633 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5192__B _5198_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_847 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3705__B _3703_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_195 VGND VPWR sky130_fd_sc_hd__decap_12
X_4459_ _4461_/A _4459_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_666 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_10 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3856__A1 data_in1[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_945 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_591 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4817__A _4817_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5058__B1 _5056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_552 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3721__A _5524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_488 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_797 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_842 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3440__B _3402_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4255__C _4255_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_503 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_480 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_856 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__A _4944_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4033__B2 _4032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5367__B key_in[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_530 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_720 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3168__A _3169_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3685__B1_N _3727_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_747 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_780 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_920 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_493 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_930 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3615__B _3570_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_964 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5533__D _3286_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5297__B1 _5325_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_463 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_528 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_720 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3847__B2 _3846_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_753 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_775 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3631__A _3579_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_477 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_609 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_650 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4165__C _4165_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_789 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4462__A _4469_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3830_ _3785_/B _3829_/X _3830_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3378__A3 _3375_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4181__B _4182_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3761_ _3749_/Y _3782_/B _3761_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_146_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3078__A _3077_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5500_ _4042_/X _3030_/A _4363_/X _5429_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2712_ _2770_/A _2711_/Y _2712_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_72_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3692_ _3671_/X _3674_/X _3692_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_5431_ _5431_/D data_out2[29] _4444_/X _5430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_127_950 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3535__B1 _3533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3806__A _3804_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2710__A _4871_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5362_ _5361_/A _5361_/B _2719_/A _5364_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_142_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_110 VGND VPWR sky130_fd_sc_hd__decap_4
X_4313_ _4312_/A _4313_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_153_290 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5443__D _5443_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_5293_ _3626_/A _5292_/X _5274_/A _5262_/X _5294_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_99_377 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_474 VGND VPWR sky130_fd_sc_hd__decap_12
X_4244_ _4244_/A _4243_/X _4244_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_99_399 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_742 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_764 VGND VPWR sky130_fd_sc_hd__decap_4
X_4175_ _4172_/X _4174_/B _4174_/X _4175_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_95_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4637__A _4637_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3541__A _3489_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_583 VGND VPWR sky130_fd_sc_hd__fill_2
X_3126_ _4985_/X _3081_/B _3129_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_458 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_778 VGND VPWR sky130_fd_sc_hd__decap_12
X_3057_ _3051_/Y _3057_/B _3055_/Y _3056_/Y _3057_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_24_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_300 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_867 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4082__A1_N _3299_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4372__A _4375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_839 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_878 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_163 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_530 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4091__B _4090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_185 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_38 VGND VPWR sky130_fd_sc_hd__decap_8
X_3959_ _3909_/X _3936_/X _3912_/Y _3959_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_149_574 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3774__B1 _3636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_769 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3716__A _3712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4869__A3 _4868_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_215 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3435__B _3432_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_655 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_986 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_699 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_720 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_742 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5545__RESET_B _4308_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4547__A _4874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_628 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5440__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_425 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_959 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_296 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3170__B _3170_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_52 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_918 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4254__A1 _4578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_789 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_85 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_694 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2804__A2 _2772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_182 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_491 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_61 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4282__A _4276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_72 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_141 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_83 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_984 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_686 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__B _5098_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5528__D _3101_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_196 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_703 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_883 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3329__C _3258_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_510 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_758 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_clock clkbuf_2_2_0_clock/X clkbuf_4_9_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_157_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_503 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3626__A _3626_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3345__B _3297_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4190__B1 _4174_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3532__A3 _3529_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_804 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_975 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4936__B1_N _4949_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_826 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_848 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_647 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4457__A _4461_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_915 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_252 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3361__A _3361_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_594 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_745 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_767 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_778 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_553 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_715 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4245__B2 _4244_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_597 VGND VPWR sky130_fd_sc_hd__decap_12
X_4931_ _4870_/X _4928_/X _4929_/Y _2907_/A _4930_/X _5458_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4796__A2 _4674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4904__B _4902_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_940 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5288__A _5288_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4862_ _4545_/A _4861_/X _4545_/A _4861_/X _4862_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__2705__A _5299_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_314 VGND VPWR sky130_fd_sc_hd__decap_12
X_3813_ _3569_/A _3835_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4793_ _3300_/A _4674_/A data_out1[28] _4677_/A _4793_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__5438__D _4643_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_714 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3756__B1 _2796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4920__A _2907_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3744_ _3743_/X _3744_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4953__C1 _4952_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_747 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_909 VGND VPWR sky130_fd_sc_hd__decap_6
X_3675_ _3674_/A _3674_/B _3675_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_106_419 VGND VPWR sky130_fd_sc_hd__fill_2
X_5414_ _5414_/D data_out2[12] _4465_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_739 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_780 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_569 VGND VPWR sky130_fd_sc_hd__decap_12
X_5345_ _2769_/A _5345_/B _5345_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_463 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_997 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5463__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_5276_ _5253_/Y _5276_/B _5276_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_336 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_196 VGND VPWR sky130_fd_sc_hd__fill_2
X_4227_ _3535_/X _4226_/X _3535_/X _4226_/X _4227_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4367__A _4367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3271__A _3270_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_937 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_414 VGND VPWR sky130_fd_sc_hd__decap_12
X_4158_ _3396_/X _4154_/X _4157_/Y _4158_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4086__B _4113_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_745 VGND VPWR sky130_fd_sc_hd__fill_1
X_3109_ _2961_/A _3108_/A _3870_/A _3108_/Y _3110_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_4089_ data_in1[23] _3976_/X _4071_/X _4088_/Y _4089_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_55_266 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3039__A2 _3037_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_737 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4814__B _4812_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4787__A2 _4781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_631 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5198__A _5198_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_642 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2798__A1 _3671_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2798__B2 _2961_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_664 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_461 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_995 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_314 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3747__B1 _3719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4830__A _4830_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_831 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_875 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_341 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5333__A1_N _5325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_257 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_717 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2988__C _2924_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4172__B1 _5534_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4711__A2 _4699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_761 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_923 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5348__A1_N _5324_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_422 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3058__A2_N _3057_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4277__A _4276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_306 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3278__A2 _3274_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_756 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4227__B2 _4226_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_981 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_480 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__B1 _3984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_483 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_157 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3738__B1 _3720_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_678 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_330 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3356__A _3356_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_514 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5486__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3460_ _3317_/X _3458_/Y _3460_/C _3460_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_143_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_867 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4702__A2 _4699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5467__RESET_B _4401_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3391_ _5222_/A _3391_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_170_377 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2713__B2 _2712_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5130_ _5052_/A _5130_/B _5130_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_69_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5290__B _5290_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4187__A _4073_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5061_ _5059_/A _5058_/X _5061_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_477 VGND VPWR sky130_fd_sc_hd__decap_8
X_4012_ _3999_/Y _4011_/X _3999_/Y _4011_/X _4012_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_531 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_704 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_406 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_258 VGND VPWR sky130_fd_sc_hd__fill_2
X_4914_ _4886_/X _4914_/B _4888_/X _4914_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_21_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_4845_ _4802_/X _4843_/Y _4844_/X _4836_/A _4815_/X _4845_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_21_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_319 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_144 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4650__A _4524_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_511 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_166 VGND VPWR sky130_fd_sc_hd__decap_8
X_4776_ _4775_/X _4769_/X data_out1[19] _4770_/X _4776_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_158_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_544 VGND VPWR sky130_fd_sc_hd__fill_1
X_3727_ _3727_/A _3704_/X _3727_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4941__A2 _4847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3266__A _5469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_588 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_845 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_396 VGND VPWR sky130_fd_sc_hd__fill_1
X_3658_ _3681_/A _3680_/A _3658_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__4154__B1 _4151_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3589_ _5517_/Q _3589_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_761 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2704__A1 _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_623 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3901__B1 _3882_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5328_ _5327_/X _5332_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_731 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_422 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4809__B _4809_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_764 VGND VPWR sky130_fd_sc_hd__fill_2
X_5259_ _3608_/A _2717_/A _5230_/X _5258_/Y _5274_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4097__A _5540_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_306 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_892 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3432__C _3432_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_767 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4825__A _4822_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_406 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_884 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4209__A1 _3980_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_417 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4209__B2 _4190_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_288 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_748 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_534 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4544__B _4542_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_940 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_422 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4263__C _4258_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_483 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_111 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_617 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_965 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_105 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4560__A _5197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5272__A1_N _5264_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2999__B _2999_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_159 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_363 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3176__A _3060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_525 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4145__B1 _4720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5560__RESET_B _4291_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_866 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_601 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_377 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3904__A _3794_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_634 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_753 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5541__D _3546_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5210__A1_N _4811_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4924__A2_N _4923_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_542 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_81 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_726 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_748 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_556 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_409 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_578 VGND VPWR sky130_fd_sc_hd__fill_2
X_2960_ _2819_/A _2959_/A _3778_/A _3158_/A _2961_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_15_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_781 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_954 VGND VPWR sky130_fd_sc_hd__fill_2
X_2891_ _2714_/Y _2891_/B _2945_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_442 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4470__A _4475_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4630_ _4630_/A _4631_/A VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_998 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5285__B _5275_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_4561_ _5562_/Q _4561_/B _4561_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2702__B _2690_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3512_ _3493_/C _3539_/B _3540_/B _3513_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3517__C _3517_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_845 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_396 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A clkbuf_3_2_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4492_ _4492_/A _4492_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_878 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_344 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4136__B1 _3382_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_569 VGND VPWR sky130_fd_sc_hd__decap_8
X_3443_ _3499_/A key_in[59] _3443_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_528 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3814__A _3793_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3374_ _3334_/X key_in[57] _3374_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4629__B _4629_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_442 VGND VPWR sky130_fd_sc_hd__fill_2
X_5113_ _5113_/A _5111_/X _5114_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_112_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5451__D _4845_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_915 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_797 VGND VPWR sky130_fd_sc_hd__decap_12
X_5044_ _5056_/A _5057_/B _5047_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_57_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_285 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_296 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3111__A1 _3110_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5501__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4645__A _4644_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_737 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_320 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3690__A1_N _3681_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_718 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_578 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_904 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_239 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_937 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_4828_ _4541_/A _4818_/X _4819_/A _4828_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_22_987 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4380__A _4381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5195__B _5192_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5389__RESET_B _4494_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4759_ _3778_/A _4757_/X data_out1[10] _4758_/X _4759_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_107_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_300 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4678__A1 _3573_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3724__A _3723_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_921 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4678__B2 _4677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2689__B1 _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_335 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_442 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3443__B key_in[59] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3350__A1 _3321_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3350__B2 _3419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4258__C _4258_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_274 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_clock clkbuf_4_3_0_clock/A _5430_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_296 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_169 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4555__A _4555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_575 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_361 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3653__A2 _3581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_707 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_898 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_217 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_220 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_792 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_903 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_431 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3810__C1 _3809_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_264 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_751 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_402 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4290__A _4304_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_436 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_297 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3618__B _3634_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5536__D _3390_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_479 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_480 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3914__B1_N _3913_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_697 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3634__A _3634_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_184 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3353__B _3356_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_453 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5524__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_924 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_328 VGND VPWR sky130_fd_sc_hd__fill_2
X_3090_ _3090_/A _3038_/X _3090_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_66_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_873 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4465__A _4468_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_501 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4841__A1 _4840_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3644__A2 _3640_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_534 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_718 VGND VPWR sky130_fd_sc_hd__fill_2
X_3992_ _4775_/X _3990_/X _4018_/B _4015_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_22_239 VGND VPWR sky130_fd_sc_hd__decap_6
X_2943_ _2943_/A _2943_/B _2944_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_31_751 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3809__A _3788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5296__A _5296_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2874_ _3801_/A _2873_/X _3801_/A _2873_/X _2887_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_918 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2805__A1_N _2814_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4613_ _5446_/Q _4610_/X _5446_/Q _4610_/X _4613_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__3528__B key_in[62] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5482__RESET_B _4384_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_661 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5446__D _4613_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_980 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5411__RESET_B _4468_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4544_ _5548_/Q _4542_/B _5548_/D VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3247__C _4720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_491 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_653 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4109__B1 _3347_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3580__A1 data_in1[0] VGND VPWR sky130_fd_sc_hd__diode_2
X_4475_ _4475_/A _4475_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_19 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3544__A _3543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_388 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_848 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_314 VGND VPWR sky130_fd_sc_hd__fill_2
X_3426_ _3361_/A _3388_/B _3359_/Y _3426_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_143_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3263__B key_in[86] VGND VPWR sky130_fd_sc_hd__diode_2
X_3357_ _3206_/X _3357_/B _3357_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_86_924 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_957 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_445 VGND VPWR sky130_fd_sc_hd__decap_6
X_3288_ _3288_/A _3285_/B _3312_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_57_158 VGND VPWR sky130_fd_sc_hd__decap_12
X_5027_ _5027_/A _5027_/B _5027_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4375__A _4375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_670 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_180 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4094__B _4093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_331 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_651 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_729 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_695 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3719__A _3765_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_272 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3438__B _3464_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_981 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4260__D _4263_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_951 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_193 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_130 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_664 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5547__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_815 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2996__C _3020_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_623 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3323__A1 _3180_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3323__B2 _3495_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_870 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_61 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4285__A _4289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_139 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_556 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_813 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_375 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_60 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3629__A _3630_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_261 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_778 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3535__A1_N _3533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_428 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4170__D _4170_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_439 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_81 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3011__B1 _3804_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_163 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3364__A _3216_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_623 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4172__A2_N _4731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_634 VGND VPWR sky130_fd_sc_hd__fill_2
X_4260_ _4616_/X _4659_/Y _4255_/C _4263_/D _4260_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_99_548 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3868__B1_N _3815_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_559 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4179__B _4177_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3314__A1 data_in2[23] VGND VPWR sky130_fd_sc_hd__diode_2
X_3211_ _3206_/X _3210_/Y _3211_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_140_166 VGND VPWR sky130_fd_sc_hd__decap_6
X_4191_ _4189_/Y _4190_/X _4191_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_39_103 VGND VPWR sky130_fd_sc_hd__decap_12
X_3142_ data_in2[18] _2956_/X _3103_/X _3141_/Y _3142_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_95_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5067__B2 _5066_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_3073_ _3026_/A _2884_/B _3073_/C _3073_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_67_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_810 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_832 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_128 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_802 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_813 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4923__A _4921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_3975_ data_in1[18] _3837_/X _3950_/X _3974_/Y _5497_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_50_345 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4042__A2 _3976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3539__A _3493_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2926_ _2925_/A _2924_/Y _2926_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_149_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_778 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3258__B _3258_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2857_ _5358_/A _2887_/A _2857_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_148_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_748 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_940 VGND VPWR sky130_fd_sc_hd__decap_8
X_5576_ _5576_/D _4524_/A _4271_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_631 VGND VPWR sky130_fd_sc_hd__decap_12
X_2788_ _5301_/A _2790_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3553__A1 _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4527_ _4577_/A _4578_/A _4525_/X _4629_/D _4527_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_172_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_4458_ _4461_/A _4458_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_105_859 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_807 VGND VPWR sky130_fd_sc_hd__fill_2
X_3409_ _3499_/A key_in[122] _3408_/X _3409_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_59_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_209 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_924 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_870 VGND VPWR sky130_fd_sc_hd__fill_2
X_4389_ _4387_/A _4389_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_570 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3856__A2 _3837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_434 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_520 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5058__A1 _5030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5058__B2 _5057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_810 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_286 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_21 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4255__D _4254_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_971 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_813 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_150 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4833__A _4833_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_515 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__B _4547_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_69 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_30 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3964__A2_N _3963_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_890 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3168__B _3169_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_918 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_732 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_703 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_597 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_758 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_769 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_601 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_675 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_995 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3184__A _3115_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_163 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_634 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3615__C _5260_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_953 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5297__A1 _5294_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_975 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1002 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_412 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3912__A _3889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_765 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_927 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3631__B _3631_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_787 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_798 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_clock clkbuf_2_0_0_clock/X clkbuf_4_1_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_65_949 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_854 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_342 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_662 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_971 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3480__B1 _3469_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_879 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3359__A _3359_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_520 VGND VPWR sky130_fd_sc_hd__decap_6
X_3760_ _3759_/A _3758_/X _3759_/X _3782_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3232__B1 _3113_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2711_ _4871_/A _2711_/B _2711_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3078__B key_in[81] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_929 VGND VPWR sky130_fd_sc_hd__decap_12
X_3691_ _4750_/X _3690_/X _4750_/X _3690_/X _3694_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5430_ _4733_/X data_out2[28] _4445_/X _5430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_65_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3806__B _3805_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3535__B2 _3534_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4732__B1 data_out2[27] VGND VPWR sky130_fd_sc_hd__diode_2
X_5361_ _5361_/A _5361_/B _2719_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2710__B _2711_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_943 VGND VPWR sky130_fd_sc_hd__decap_3
X_4312_ _4312_/A _4312_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5292_ _5262_/B _5292_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_367 VGND VPWR sky130_fd_sc_hd__decap_3
X_4243_ _4241_/X _4242_/X _4243_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__4918__A _4918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3299__B1 _3297_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3822__A _3818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_188 VGND VPWR sky130_fd_sc_hd__fill_2
X_4174_ _4172_/X _4174_/B _4174_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3541__B _3513_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3125_ _4996_/A _3122_/X _3124_/Y _3125_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_95_573 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_938 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_798 VGND VPWR sky130_fd_sc_hd__fill_2
X_3056_ _2911_/X _3055_/B _3056_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_35_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_982 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4653__A _4577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_429 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_790 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5212__A1 _5211_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5392__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_328 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_507 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3269__A _3228_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_378 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_389 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3223__B1 _3222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_542 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4091__C _4786_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3958_ _3133_/A _3956_/X _3957_/X _3958_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3774__A1 _3724_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1007 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3774__B2 _3751_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2909_ _2838_/A _2865_/X _2836_/Y _2909_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_137_726 VGND VPWR sky130_fd_sc_hd__decap_6
X_3889_ _3770_/Y _3887_/X _3889_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_109_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_718 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3716__B _3714_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4723__B1 data_out2[23] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_589 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_910 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_984 VGND VPWR sky130_fd_sc_hd__decap_4
X_5559_ _5559_/D _4997_/C _4292_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_118_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_227 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_177 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3732__A _3661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_754 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4547__B _4547_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_873 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_949 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3170__C _3170_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_64 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_802 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_971 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_407 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4254__A2 _4252_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_97 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4563__A _5564_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5514__RESET_B _4345_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_930 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_879 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_73 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_816 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_339 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_95 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_849 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_715 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_737 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3907__A _3062_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_50 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_573 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_556 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_718 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_578 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3626__B _3625_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4714__B1 data_out2[18] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5544__D _4540_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_228 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_483 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4190__A1 _3955_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3345__C _3271_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_261 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3642__A _3641_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_702 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_562 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3361__B _3359_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_448 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_908 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_407 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4473__A _4475_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4930_ _4815_/A _4930_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3453__B1 _3442_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_952 VGND VPWR sky130_fd_sc_hd__decap_12
X_4861_ _5548_/Q _4849_/X _4873_/A _4861_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_61_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2705__B key_in[39] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_687 VGND VPWR sky130_fd_sc_hd__decap_12
X_3812_ _3765_/A _3812_/B _2714_/A _3812_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4792_ _4791_/X _4781_/X data_out1[27] _4782_/X _4792_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_20_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3756__B2 _3755_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3743_ _3740_/X _3742_/X _3743_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4953__B1 _4942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_726 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_895 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3817__A _2918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_737 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_545 VGND VPWR sky130_fd_sc_hd__fill_1
X_3674_ _3674_/A _3674_/B _3674_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3508__A1 _3505_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5413_ _5413_/D data_out2[11] _4466_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5454__D _4881_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_537 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_792 VGND VPWR sky130_fd_sc_hd__fill_1
X_5344_ _5343_/X _5345_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_773 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3351__A1_N _3316_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_261 VGND VPWR sky130_fd_sc_hd__fill_2
X_5275_ _5256_/Y _5275_/B _5276_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__4648__A _4645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_626 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3552__A _3529_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4226_ _4225_/A _4224_/X _4225_/X _4226_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_29_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_871 VGND VPWR sky130_fd_sc_hd__decap_12
X_4157_ _4156_/X _4157_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_28_426 VGND VPWR sky130_fd_sc_hd__decap_12
X_3108_ _3108_/A _3108_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_28_459 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_554 VGND VPWR sky130_fd_sc_hd__decap_8
X_4088_ _3974_/A _4088_/B _4087_/X _4088_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_83_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_576 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_278 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4383__A _4397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_289 VGND VPWR sky130_fd_sc_hd__fill_2
X_3039_ _3038_/A _3037_/Y _3038_/X _3039_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_70_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_56 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5198__B _5198_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_16 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2798__A2 _3870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_626 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_676 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_125 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3747__A1 data_in1[8] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4830__B _4830_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2955__C1 _2954_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3727__A _3727_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_31 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4172__B2 _5538_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_827 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_464 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4558__A _4987_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3462__A _3519_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_540 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_702 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_871 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_882 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_74 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3683__B1 _5513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_381 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4293__A _4296_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2806__A _2847_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_749 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_952 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3986__B2 _3985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5539__D _5539_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_760 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_771 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_613 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_136 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_624 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5188__B1 _5185_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_495 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3738__B2 _3737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_821 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_842 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_875 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3356__B _3356_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5360__B1 _5481_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_879 VGND VPWR sky130_fd_sc_hd__decap_12
X_3390_ data_in2[25] _3172_/X _3364_/X _3389_/Y _3390_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_170_389 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4468__A _4468_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_570 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3165__A2_N _3164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4081__A1_N _4079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_592 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3372__A _3326_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5060_ _5072_/B _5060_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_85_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_979 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4187__B _4187_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4011_ _3200_/X _4010_/X _3200_/X _4010_/X _4011_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5436__RESET_B _4438_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_223 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_234 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_768 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_351 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5299__A _5299_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_598 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2716__A _2716_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_481 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_557 VGND VPWR sky130_fd_sc_hd__fill_2
X_4913_ _4900_/A _4899_/X _4885_/Y _4913_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__5449__D _4826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_760 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_782 VGND VPWR sky130_fd_sc_hd__fill_2
X_4844_ _4841_/X _4842_/X _4844_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_635 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_629 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_668 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4650__B _4650_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_681 VGND VPWR sky130_fd_sc_hd__fill_2
X_4775_ _2959_/A _4775_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3726_ _2735_/X _3722_/X _3725_/Y _3726_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__4034__A1_N _3230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5430__CLK _5430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3266__B _3266_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_729 VGND VPWR sky130_fd_sc_hd__decap_3
X_3657_ _3634_/X _3657_/B _3680_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_857 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4154__B2 _4153_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3588_ _3588_/A _3588_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_161_367 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2704__A2 _2688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3901__A1 data_in1[15] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4378__A _4381_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5327_ _5327_/A _5327_/B _5327_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_142_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_743 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_123 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5103__B1 _5569_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_5258_ _5258_/A _5258_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4209_ _3980_/Y _3463_/Y _4188_/X _4190_/X _4209_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_5189_ _4798_/B _5189_/B _5211_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_29_757 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4825__B _4825_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4209__A2 _3463_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_429 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_790 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5002__A _5001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_974 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4263__D _4263_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_270 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_495 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_617 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_679 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_999 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2928__C1 _2927_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3457__A _3488_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_138 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_898 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3176__B _3176_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_684 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_375 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_323 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_397 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_183 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_322 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4145__A1 _3932_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4145__B2 _3548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1000 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_507 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3904__B _3903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_388 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4288__A _4289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_646 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_819 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_253 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3920__A _3872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_61 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_259 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4081__B1 _4079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_473 VGND VPWR sky130_fd_sc_hd__fill_2
X_2890_ _5292_/X _2889_/A _5261_/A _2889_/Y _2891_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__5453__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_977 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_821 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_320 VGND VPWR sky130_fd_sc_hd__decap_12
X_4560_ _5197_/A _4561_/B VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_301 VGND VPWR sky130_fd_sc_hd__decap_4
X_3511_ _3493_/C _3539_/B _3540_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4491_ _4492_/A _4491_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_7_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4136__B2 _4135_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3442_ _3441_/A _3441_/B _3441_/X _3442_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_6_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5333__B1 _5325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_922 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3814__B _3802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4198__A _4198_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3373_ _3371_/X _3372_/X _3371_/X _3372_/X _3373_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4629__C _4578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_220 VGND VPWR sky130_fd_sc_hd__fill_2
X_5112_ _5113_/A _5111_/X _5114_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_69_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_476 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_253 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_776 VGND VPWR sky130_fd_sc_hd__decap_6
X_5043_ _5036_/Y _5040_/X _5057_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_69_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_938 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_498 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3830__A _3785_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_137 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3111__A2 _3110_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_822 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_693 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_749 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_332 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4661__A _5198_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_933 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_793 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_607 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5347__A1_N _5333_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_955 VGND VPWR sky130_fd_sc_hd__decap_3
X_4827_ _4827_/A _4830_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_138_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3277__A _3288_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_448 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5195__C _5194_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4758_ _4701_/A _4758_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_1000 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_802 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_515 VGND VPWR sky130_fd_sc_hd__decap_8
X_3709_ _2713_/X _3708_/X _2713_/X _3708_/X _3709_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_621 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_312 VGND VPWR sky130_fd_sc_hd__fill_2
X_4689_ _5356_/C _4687_/X data_out2[6] _4688_/X _4689_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_162_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_183 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_507 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4678__A2 _4674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_721 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2689__B2 _2688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3886__B1 _3860_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_955 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3350__A2 _3349_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_819 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_476 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_787 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_627 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4836__A _4836_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_47 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4555__B _4541_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_52 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_844 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5476__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_771 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_782 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_221 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4571__A _5571_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_232 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3810__B1 _3790_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_265 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_977 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_276 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_62 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5012__C1 _5011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_84 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3187__A _3187_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_971 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_643 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_631 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4812__B1_N _4823_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_378 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3634__B _3624_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5552__D _4549_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5131__A2_N _5130_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_402 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_318 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4746__A _4701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_881 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3650__A _3651_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_608 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4841__A2 _4839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_3991_ _4775_/X _3990_/X _4018_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5251__C1 _5250_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_771 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4481__A _4477_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_549 VGND VPWR sky130_fd_sc_hd__fill_1
X_2942_ _2943_/A _2943_/B _2944_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_95_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_916 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3809__B _3807_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_949 VGND VPWR sky130_fd_sc_hd__decap_12
X_2873_ _2871_/X _2872_/X _2871_/X _2872_/X _2873_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_4612_ _4646_/B _4609_/B _4611_/Y _4612_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_157_982 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_150 VGND VPWR sky130_fd_sc_hd__decap_3
X_4543_ _5547_/Q _4542_/B _5547_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_129_695 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5306__B1 _4836_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4109__B2 _4108_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_974 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_665 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_805 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3580__A2 _3391_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4474_ _4475_/A _4474_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3544__B _3543_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5451__RESET_B _4421_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3425_ _3395_/X _3421_/X _3435_/A _3431_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__5462__D _5462_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3356_ _3356_/A _3356_/B _3357_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_947 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_830 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4656__A _4655_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3287_ _3216_/A _3143_/B _3287_/C _3287_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5499__CLK _5430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_5026_ _5563_/Q _5025_/X _5563_/Q _5025_/X _5027_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_800 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_362 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_129 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_844 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_343 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4391__A _4390_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_538 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2904__A _2904_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_201 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3719__B _3679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_223 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_757 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_971 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_918 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_835 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_621 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_428 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5539__RESET_B _4315_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_54 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_323 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3735__A _3734_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_98 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_827 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_623 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5372__D _4743_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3859__B1 _2842_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_741 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3323__A2 _3322_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_763 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_627 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_936 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4566__A _4566_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_435 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5239__A1_N _4817_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3470__A _3499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_479 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_928 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_991 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_877 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_579 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_888 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4036__B1 _4034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2814__A _2702_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_858 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_701 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3629__B _3628_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_763 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5547__D _5547_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_960 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_407 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_470 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3011__A1 _2870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3011__B2 _3180_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_816 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3364__B _3364_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2773__A2_N _2772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_657 VGND VPWR sky130_fd_sc_hd__fill_2
X_3210_ _3207_/X _3210_/B _3209_/Y _3210_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_5_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3314__A2 _3172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_679 VGND VPWR sky130_fd_sc_hd__fill_2
X_4190_ _3955_/Y _4047_/Y _4174_/X _4190_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3141_ _3170_/A _3139_/Y _3141_/C _3141_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_39_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_947 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4476__A _4469_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_733 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_766 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_243 VGND VPWR sky130_fd_sc_hd__decap_12
X_3072_ data_in2[16] _2956_/X _3026_/X _3071_/Y _5527_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_83_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_660 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4923__B _4922_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_162 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_538 VGND VPWR sky130_fd_sc_hd__decap_8
X_3974_ _3974_/A _3972_/Y _3973_/X _3974_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__5100__A _5473_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_724 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3539__B _3539_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2925_ _2925_/A _2924_/Y _2925_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5457__D _4919_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_757 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3258__C _3258_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2856_ _2814_/X _2840_/X _2887_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_108_109 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_237 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_790 VGND VPWR sky130_fd_sc_hd__decap_3
X_5575_ _4255_/X _4650_/B _4272_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2787_ _2898_/A key_in[41] _2787_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_643 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3553__A2 key_in[127] VGND VPWR sky130_fd_sc_hd__diode_2
X_4526_ _4650_/B _4629_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_827 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_4457_ _4461_/A _4457_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_3408_ _3222_/X _3408_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_167 VGND VPWR sky130_fd_sc_hd__fill_2
X_4388_ _4387_/A _4388_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3339_ _4639_/X _3335_/X _3336_/X _3337_/X _3338_/X _3340_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_59_958 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4386__A _4387_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_381 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3290__A _4582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5058__A2 _5047_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_265 VGND VPWR sky130_fd_sc_hd__decap_8
X_5009_ _5008_/X _5009_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_298 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_983 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4833__B _4833_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_162 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_994 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_387 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_549 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_99 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5010__A _5009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_20 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5514__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4862__A2_N _4861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_744 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_755 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_418 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_226 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2866__A1_N _2858_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5373__RESET_B _4513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_236 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3465__A _3465_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_131 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_462 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3184__B _3185_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_977 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5297__A2 _5294_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_307 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_571 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3912__B _3910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_582 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_733 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2809__A _2784_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4296__A _4296_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3631__C _3630_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_619 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_800 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4257__B1 _4256_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_939 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_747 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_310 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2807__A1 _2847_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_641 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_961 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_814 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3480__B2 _3479_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_666 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3359__B _3359_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3232__A1 _2889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_571 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3232__B2 _3231_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_70 VGND VPWR sky130_fd_sc_hd__decap_3
X_2710_ _4871_/A _2711_/B _2770_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_158_565 VGND VPWR sky130_fd_sc_hd__decap_12
X_3690_ _3681_/Y _3689_/Y _3681_/Y _3689_/Y _3690_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_941 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3375__A _3337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4732__A1 _4731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_974 VGND VPWR sky130_fd_sc_hd__fill_2
X_5360_ _3608_/A _3804_/A _5481_/Q _2870_/A _5361_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_127_985 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4732__B2 _4726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_770 VGND VPWR sky130_fd_sc_hd__fill_2
X_4311_ _4304_/A _4312_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_421 VGND VPWR sky130_fd_sc_hd__fill_2
X_5291_ _5290_/A _5290_/B _5325_/A _5294_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_114_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_454 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_519 VGND VPWR sky130_fd_sc_hd__decap_4
X_4242_ _4047_/Y _5542_/Q _4731_/X _3548_/Y _4242_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4918__B _4916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3299__B2 _3298_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_178 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3822__B _3821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4173_ _4146_/X _4173_/B _4174_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_110_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2719__A _2719_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_541 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_777 VGND VPWR sky130_fd_sc_hd__fill_2
X_3124_ _3124_/A _3124_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3541__C _3541_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4248__B1 data_in1[31] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_3055_ _2910_/Y _3055_/B _3055_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_48_490 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_909 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_825 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_994 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4653__B _4522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_696 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5537__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_324 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_357 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5212__A2 _5210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3269__B _3226_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_519 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3223__A1 _3291_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3957_ _3133_/A _3956_/X _3957_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_18 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3774__A2 _3752_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2908_ _2832_/A _2864_/X _2908_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_390 VGND VPWR sky130_fd_sc_hd__fill_2
X_3888_ _3770_/Y _3887_/X _3888_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_13_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_2839_ _2838_/A _2837_/X _2838_/X _2839_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3285__A _3170_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4184__C1 _4183_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4723__A1 _3287_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_5558_ _4555_/X _4555_/A _4293_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4723__B2 _4713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_4509_ _4504_/X _4509_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_105_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_292 VGND VPWR sky130_fd_sc_hd__decap_12
X_5489_ _3789_/X _4756_/A _4375_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_133_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_796 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3732__B _3730_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_830 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_766 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5005__A _4982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_863 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_574 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4239__B1 _3397_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_276 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3852__B1_N _3851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_747 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4844__A _4841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_630 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_652 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4563__B _4557_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_994 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_324 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_52 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_290 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_357 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_368 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5554__RESET_B _4298_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_841 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_176 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_204 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_384 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_535 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3907__B _3906_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_941 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3195__A _5013_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_952 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4714__A1 _5529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4714__B2 _4713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_410 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_281 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_421 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4190__A2 _4047_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_292 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3923__A _3874_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_349 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5560__D _5560_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3150__B1 _3148_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5040__A1_N _5564_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_939 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4754__A _5288_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_611 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3453__B2 _3452_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_4860_ _4819_/A _4873_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_644 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_964 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_3811_ _4664_/X _3812_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_4791_ _3251_/A _4791_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_699 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_187 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_390 VGND VPWR sky130_fd_sc_hd__decap_8
X_3742_ _2717_/A _3710_/X _3741_/X _3742_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__4953__A1 _4943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3817__B _3816_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_383 VGND VPWR sky130_fd_sc_hd__decap_8
X_3673_ _3647_/X _3651_/X _3674_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_5412_ _4695_/X data_out2[10] _4467_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3508__A2 _3507_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4166__C1 _4165_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_760 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_410 VGND VPWR sky130_fd_sc_hd__fill_2
X_5343_ _5342_/X _5343_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4929__A _4928_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3833__A _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_839 VGND VPWR sky130_fd_sc_hd__decap_4
X_5274_ _5274_/A _5274_/B _5275_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_130_936 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_104 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_947 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3552__B key_in[95] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_295 VGND VPWR sky130_fd_sc_hd__fill_2
X_4225_ _4225_/A _4224_/X _4225_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5470__D _5075_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_703 VGND VPWR sky130_fd_sc_hd__decap_4
X_4156_ _4155_/X _4156_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_95_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_725 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_736 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_438 VGND VPWR sky130_fd_sc_hd__decap_12
X_3107_ _3060_/A _3107_/B _3107_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4664__A _3584_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4087_ _4072_/Y _4113_/B _4087_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3348__A2_N _3347_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_961 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_408 VGND VPWR sky130_fd_sc_hd__decap_12
X_3038_ _3038_/A _3037_/Y _3038_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4641__B1 _5448_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_791 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_121 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_688 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_839 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4989_ _4985_/X _4987_/X _4988_/X _4992_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2912__A _2910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3747__A2 _3697_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_861 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2955__B1 _2929_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3727__B _3704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_855 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_43 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4839__A _5547_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_741 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_559 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3743__A _3740_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4558__B _4557_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_593 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_284 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3462__B _3364_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5380__D _4759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3132__B1 _3107_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_660 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3683__A1 _3603_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_894 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3683__B2 _3682_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4574__A _5165_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_717 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2806__B _2847_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_791 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_964 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_666 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A1 _4635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_783 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5188__B2 _5187_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_636 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3918__A _3032_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2822__A _2822_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3411__A1_N _5473_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_693 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_61 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_872 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2946__B1 _2964_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_894 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5555__D _4552_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_505 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_527 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_324 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5360__A1 _3608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5360__B2 _2870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3372__B _3331_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5382__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_338 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_2_0_clock_A clkbuf_4_3_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_4010_ _4003_/X _4008_/Y _4009_/X _4010_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_77_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_980 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4484__A _4483_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2882__C1 _2881_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_961 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_257 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_363 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5476__RESET_B _4391_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2716__B _2717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_238 VGND VPWR sky130_fd_sc_hd__fill_2
X_4912_ _4911_/A _4910_/X _4911_/X _4917_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_18_493 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5405__RESET_B _4475_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_441 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_772 VGND VPWR sky130_fd_sc_hd__decap_8
X_4843_ _4841_/X _4842_/X _4843_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_61_794 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3828__A _3828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2732__A _5223_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4926__A1 _4925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_658 VGND VPWR sky130_fd_sc_hd__decap_4
X_4774_ _5497_/Q _4769_/X data_out1[18] _4770_/X _4774_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_147_822 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4650__C _4518_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3725_ _3724_/X _3725_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_20_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_855 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5465__D _5012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_814 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_825 VGND VPWR sky130_fd_sc_hd__decap_4
X_3656_ _3645_/X _3657_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_869 VGND VPWR sky130_fd_sc_hd__decap_12
X_3587_ _3575_/X _3587_/B _3587_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3272__A2_N _3271_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_5326_ _5199_/Y _4756_/A _5199_/Y _4756_/A _5327_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_774 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3901__A2 _3837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_755 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5103__B2 _5102_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5257_ _2716_/A _2717_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3114__B1 _3113_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_319 VGND VPWR sky130_fd_sc_hd__decap_12
X_4208_ _4728_/X _3493_/C _4207_/X _4208_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_102_479 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_5188_ _4635_/A _5183_/X _5184_/X _5185_/X _5187_/X _5189_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4862__B1 _4545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_12 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2907__A _2907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4394__A _4390_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4139_ _4788_/X _4137_/X _4138_/X _4159_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_113_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_864 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_886 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3417__A1 _3416_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_739 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_558 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_964 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_614 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_102 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_945 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_282 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_800 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_629 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_822 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2928__B1 _2884_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3457__B _3457_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_844 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5375__D _5375_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_64 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3176__C _3162_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_53 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_516 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_195 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4145__A2 _5542_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4569__A _5569_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_741 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1012 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_356 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_560 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_378 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_796 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_658 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_766 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_500 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_831 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3920__B _3896_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2817__A _5494_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_834 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_441 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_761 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4081__B2 _4080_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_967 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_293 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4109__A1_N _3347_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_118 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2919__B1 _2930_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_129 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_488 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_855 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_332 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_803 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3592__B1 _5213_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3510_ _3510_/A _3510_/B _3539_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_155_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_376 VGND VPWR sky130_fd_sc_hd__decap_12
X_4490_ _4269_/A _4492_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_128_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_869 VGND VPWR sky130_fd_sc_hd__fill_2
X_3441_ _3441_/A _3441_/B _3441_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4479__A _4477_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5333__B2 _5332_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3372_ _3326_/Y _3331_/X _3372_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_934 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4198__B _4198_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_198 VGND VPWR sky130_fd_sc_hd__decap_12
X_5111_ _5086_/Y _5108_/X _5110_/X _5111_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4629__D _4629_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_135 VGND VPWR sky130_fd_sc_hd__decap_8
X_5042_ _5041_/X _5056_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_639 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3830__B _3829_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2727__A _2728_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_503 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_672 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_867 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_290 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4942__A _4546_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_878 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_772 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_591 VGND VPWR sky130_fd_sc_hd__fill_2
X_4826_ _4802_/X _4824_/Y _4832_/B _4817_/A _4815_/X _4826_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_166_427 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2892__B1_N _2945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_630 VGND VPWR sky130_fd_sc_hd__fill_2
X_4757_ _4699_/A _4757_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3708_ _3706_/X _3707_/X _3706_/X _3707_/X _3708_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4688_ _4677_/A _4688_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_173 VGND VPWR sky130_fd_sc_hd__fill_2
X_3639_ _5284_/Y _3638_/B _3666_/A _3641_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4389__A _4387_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_666 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3293__A _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_45 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3886__A1 _3861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_304 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_422 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_733 VGND VPWR sky130_fd_sc_hd__fill_2
X_5309_ _5306_/Y _5308_/X _5309_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5398__RESET_B _4484_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4835__B1 _4827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_691 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_533 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_842 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5013__A _5013_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_503 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_812 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_374 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_536 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_856 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_333 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4852__A _4852_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_86 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_200 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_377 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_794 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4571__B _4574_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3810__A1 data_in1[11] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_233 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5012__B1 _4942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_288 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_415 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_299 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3187__B _3186_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_797 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_85 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3574__B1 _3573_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_610 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5315__A1 _5284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4299__A _4303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_869 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_142 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_904 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_541 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5079__B1 _4566_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3931__A _3908_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_477 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_893 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4826__B1 _4817_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3650__B _3649_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_801 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5420__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4033__A1_N _4031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_620 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_845 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_878 VGND VPWR sky130_fd_sc_hd__fill_2
X_3990_ _3987_/X _3989_/Y _3987_/X _3989_/Y _3990_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5251__B1 _5224_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_366 VGND VPWR sky130_fd_sc_hd__fill_2
X_2941_ _2799_/A _5497_/Q _3759_/A _3110_/A _2943_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__5570__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3809__C _3808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_241 VGND VPWR sky130_fd_sc_hd__decap_4
X_2872_ _2872_/A _2822_/X _2872_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__5003__B1 _5002_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_263 VGND VPWR sky130_fd_sc_hd__fill_2
X_4611_ _4610_/X _4611_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_803 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3565__B1 _5281_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4542_ _4542_/A _4542_/B _4542_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_971 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_470 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_110 VGND VPWR sky130_fd_sc_hd__fill_2
X_4473_ _4475_/A _4473_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5306__B2 _5334_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_986 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_677 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_208 VGND VPWR sky130_fd_sc_hd__decap_6
X_3424_ _3484_/A _3435_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4002__A _3175_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3868__A1 _3794_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_3355_ _3287_/C _3309_/B _3354_/X _3359_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_112_541 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4937__A _4925_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_274 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5491__RESET_B _4373_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_736 VGND VPWR sky130_fd_sc_hd__fill_1
X_3286_ data_in2[22] _3172_/X _3247_/X _3285_/Y _3286_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_39_842 VGND VPWR sky130_fd_sc_hd__decap_12
X_5025_ _4975_/X _5024_/X _5025_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_458 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_609 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5420__RESET_B _4458_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_867 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4672__A _4671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_355 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3288__A _3288_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3719__C _5261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_235 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_909 VGND VPWR sky130_fd_sc_hd__decap_6
X_4809_ _4799_/Y _4809_/B _4810_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_11 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2920__A _2844_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_942 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_644 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_806 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3308__B1 _3290_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__A _5008_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3825__A1_N _3815_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3859__A1 _3769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5579__RESET_B _4266_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_21 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3859__B2 _3858_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_669 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_753 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4847__A _4891_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5508__RESET_B _4352_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_786 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5443__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_639 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_948 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_47 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4566__B _4561_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3470__B key_in[60] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_650 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_75 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_396 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_845 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3492__C1 _3491_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4582__A _2999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_141 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4036__B2 _4035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5233__B1 _5231_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_528 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2814__B _2722_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3198__A _3195_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_196 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3795__B1 _3819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_775 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_550 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_972 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3926__A _3925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_419 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_267 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3547__B1 _3545_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_994 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3011__A2 _3010_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_493 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_290 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_952 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5563__D _4562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_963 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_986 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_997 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3364__C _4728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_996 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_70 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_230 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4757__A _4699_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_701 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3661__A _3660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_926 VGND VPWR sky130_fd_sc_hd__decap_4
X_3140_ _3139_/A _3138_/X _3141_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__5346__A1_N _5335_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3071_ _2927_/A _3071_/B _3071_/C _3071_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_55_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_778 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_91 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4492__A _4492_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_984 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_517 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_995 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_3973_ _3972_/A _3971_/X _3973_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_51_859 VGND VPWR sky130_fd_sc_hd__fill_2
X_2924_ _2878_/A _2920_/Y _2924_/C _2923_/Y _2924_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_31_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_2855_ _2855_/A _2855_/B _2855_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_31_594 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3538__B1 _3521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_460 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2740__A _2740_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5574_ _4574_/X _5165_/A _4273_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_482 VGND VPWR sky130_fd_sc_hd__decap_6
X_2786_ _5300_/A _2898_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4525_ _4524_/Y _4525_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5473__D _5115_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_655 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_912 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_677 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3009__A2_N _3008_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_474 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5466__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_485 VGND VPWR sky130_fd_sc_hd__decap_4
X_4456_ _4461_/A _4456_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_132_625 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_349 VGND VPWR sky130_fd_sc_hd__fill_2
X_3407_ _3334_/X _3499_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4667__A _4666_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4387_ _4387_/A _4387_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3571__A _3676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_179 VGND VPWR sky130_fd_sc_hd__decap_4
X_3338_ _3334_/X key_in[120] _3222_/X _3338_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_98_594 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_222 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3290__B _3318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5058__A3 _5032_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_544 VGND VPWR sky130_fd_sc_hd__decap_8
X_3269_ _3228_/X _3226_/X _3199_/Y _3269_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_100_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5008_ _5008_/A _5006_/Y _5008_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_26_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_642 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_804 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2915__A _2915_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5215__B1 _5198_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_675 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_472 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_38 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3777__B1 _3768_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_522 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_235 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_279 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3746__A _3788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_931 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_238 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3465__B _3465_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_709 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5383__D _4764_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5145__A2_N _5144_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_923 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_466 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4577__A _4577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_403 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_319 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3912__C _3912_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_723 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_594 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2809__B _2846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_907 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_406 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4257__A1 _4517_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_288 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2807__A2 _2847_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_940 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_759 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2825__A _2934_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_686 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_612 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_483 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5558__D _4555_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_678 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3359__C _3357_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3232__A2 _3231_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_909 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_554 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_577 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3656__A _3645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5489__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_249 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4193__B1 _4187_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3375__B key_in[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_441 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4732__A2 _4725_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4310_ _4305_/A _4310_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3940__B1 _3916_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_411 VGND VPWR sky130_fd_sc_hd__decap_8
X_5290_ _5290_/A _5290_/B _5325_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_153_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_658 VGND VPWR sky130_fd_sc_hd__decap_12
X_4241_ _3395_/X _3521_/X _4225_/X _4241_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4487__A _4483_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_146 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3391__A _5222_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4918__C _4917_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4999__A2_N _4998_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4172_ _3287_/C _4731_/X _5534_/Q _5538_/Q _4172_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__2719__B _5364_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_842 VGND VPWR sky130_fd_sc_hd__decap_12
X_3123_ _4996_/A _3122_/X _3124_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_96_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_918 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4248__A1 _5197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4248__B2 _4546_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_3054_ _2975_/X _3050_/X _3055_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_36_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2735__A _2734_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_450 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_770 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_859 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_196 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5468__D _5048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3269__C _3199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4950__A _4951_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3956_ _3750_/Y _5534_/Q _2984_/A _3955_/Y _3956_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_149_522 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3223__A2 key_in[117] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3563__A2_N _3562_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2907_ _2907_/A _2863_/X _2907_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3774__A3 _3735_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3887_ _3682_/Y _3175_/A _2876_/A _3175_/Y _3887_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2982__A1 _2999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_525 VGND VPWR sky130_fd_sc_hd__decap_12
X_2838_ _2838_/A _2837_/X _2838_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_136_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3285__B _3285_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4184__B1 _4167_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5557_ _4554_/X _4554_/A _4294_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4723__A2 _4712_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2769_ _2769_/A _2767_/A _5310_/Y _2769_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_117_452 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_719 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clock_A clock VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_207 VGND VPWR sky130_fd_sc_hd__decap_3
X_4508_ _4504_/X _4508_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_794 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_422 VGND VPWR sky130_fd_sc_hd__decap_12
X_5488_ _5488_/D _5288_/A _4377_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_647 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_764 VGND VPWR sky130_fd_sc_hd__decap_8
X_4439_ _4438_/A _4439_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4397__A _4397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_775 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_606 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_56 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3732__C _3642_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_842 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5005__B _4992_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_778 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_715 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4239__B2 _3556_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_897 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4844__B _4842_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_951 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_984 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_910 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_826 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5021__A _5021_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_921 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_31 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2772__A2_N _2771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5378__D _4753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_133 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4860__A _4819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_86 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_97 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_886 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_553 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_525 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_524 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_74 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3195__B _3195_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_430 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5523__RESET_B _4335_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4714__A2 _4712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2725__A1 _5356_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_956 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_753 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3923__B _3922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_818 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2_0_clock_A clkbuf_3_2_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4100__A _4099_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3150__A1 _4638_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3150__B2 _3149_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_586 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_534 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3989__B1 _3953_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_675 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_461 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_656 VGND VPWR sky130_fd_sc_hd__fill_2
X_3810_ data_in1[11] _3697_/X _3790_/X _3809_/Y _3810_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_21_818 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4770__A _4700_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_4790_ _3231_/A _4781_/X data_out1[26] _4782_/X _4790_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_32_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_475 VGND VPWR sky130_fd_sc_hd__decap_12
X_3741_ _3741_/A _3713_/X _3741_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4953__A2 _4847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3672_ _3671_/A _3670_/X _3671_/X _3674_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_118_227 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_395 VGND VPWR sky130_fd_sc_hd__fill_2
X_5411_ _5411_/D data_out2[9] _4468_/X _5402_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4166__B1 _4144_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_772 VGND VPWR sky130_fd_sc_hd__decap_8
X_5342_ _4848_/A _5341_/B _5342_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_127_794 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4929__B _4927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3833__B _3832_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5115__C1 _5114_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_764 VGND VPWR sky130_fd_sc_hd__fill_2
X_5273_ _5263_/X _5272_/Y _5263_/X _5272_/Y _5274_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_829 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_606 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_926 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_797 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5106__A _5134_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_488 VGND VPWR sky130_fd_sc_hd__decap_12
X_4224_ _4000_/Y _4097_/Y _4207_/X _4209_/X _4224_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_99_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3677__C1 _3676_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_907 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5504__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4155_ _3396_/X _4154_/X _4155_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4945__A _4921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_512 VGND VPWR sky130_fd_sc_hd__fill_2
X_3106_ _3060_/B _3176_/B _2999_/A _3107_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_83_523 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_534 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_694 VGND VPWR sky130_fd_sc_hd__decap_8
X_4086_ _4072_/Y _4113_/B _4088_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_83_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_940 VGND VPWR sky130_fd_sc_hd__fill_2
X_3037_ _3014_/B _3037_/B _3036_/Y _3037_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_52_910 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4641__A1 _4640_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_483 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4641__B2 _4631_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_291 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_177 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4988_ _4985_/X _4987_/X _4988_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2912__B _2911_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3939_ _3794_/A _3939_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3296__A _5470_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2955__A1 data_in2[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_396 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_895 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_867 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2803__A1_N _2796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_249 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_878 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_355 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5354__C1 _5353_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_366 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_516 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_400 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_783 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_934 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4839__B _4838_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_433 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3380__A1 _5472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3743__B _3742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3462__C _5539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_531 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4829__A2_N _4828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3132__B2 _3163_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4855__A _4853_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3683__A2 _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_586 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_534 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4574__B _4574_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_951 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1009 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_729 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_740 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4590__A _4590_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_127 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A2 _5183_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3918__B _3917_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2822__B _2821_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_300 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_73 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2946__B2 _2945_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_361 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4148__B1 _4000_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3934__A _3933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_539 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_398 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5360__A2 _3804_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3371__A1 _3178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5527__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5571__D _4571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_309 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4765__A _2797_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_534 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_394 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_6_0_clock_A clkbuf_4_7_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2882__B1 _2854_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_887 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_228 VGND VPWR sky130_fd_sc_hd__fill_2
X_4911_ _4911_/A _4910_/X _4911_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_45_280 VGND VPWR sky130_fd_sc_hd__decap_12
X_4842_ _4830_/X _4842_/B _4842_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_609 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3828__B _3805_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4926__A2 _4924_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4773_ _3113_/A _4769_/X data_out1[17] _4770_/X _4773_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_165_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_136 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5445__RESET_B _4428_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_503 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4650__D _4649_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_514 VGND VPWR sky130_fd_sc_hd__fill_2
X_3724_ _3723_/X _3724_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4005__A _3958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_536 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_889 VGND VPWR sky130_fd_sc_hd__fill_1
X_3655_ _3586_/A _3681_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3533__A1_N _5154_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3844__A _3842_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_837 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_325 VGND VPWR sky130_fd_sc_hd__decap_12
X_3586_ _3586_/A _3587_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_753 VGND VPWR sky130_fd_sc_hd__decap_8
X_5325_ _5325_/A _5325_/B _5325_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_88_604 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5481__D _3614_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_572 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_712 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_5256_ _5256_/A _5256_/B _5256_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_87_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_447 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3114__A1 _3033_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4207_ _4000_/Y _4097_/Y _4207_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4675__A _4672_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5187_ _5203_/A key_in[96] _5207_/A _5187_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_68_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_981 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4862__B2 _4861_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4138_ _4788_/X _4137_/X _4138_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2907__B _2863_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2873__B1 _2871_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_57 VGND VPWR sky130_fd_sc_hd__decap_4
X_4069_ _3974_/A _4069_/B _4069_/C _4069_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3417__A2 _3415_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_39 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_431 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_902 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_436 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2923__A _2849_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_637 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_957 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_294 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2928__A1 data_in2[12] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_300 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_193 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_333 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_664 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_141 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_355 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3176__D _3163_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_65 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_697 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3754__A _3725_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_859 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4569__B _4574_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5391__D _4779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_572 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_42 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_594 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_285 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_97 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_778 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4585__A _4650_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_629 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4853__A1 _4852_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_512 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_288 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_394 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_843 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_943 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3929__A _3839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_946 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_592 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_801 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5566__D _5566_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2919__A1 _2918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_300 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_834 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_670 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_642 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_867 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3592__B2 _3591_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_837 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3664__A _3663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_314 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_388 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3347__A2_N _3346_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3440_ _3399_/X _3402_/X _3441_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_155_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_3371_ _3178_/Y _3369_/X _3370_/X _3371_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_112_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_572 VGND VPWR sky130_fd_sc_hd__fill_2
X_5110_ _5090_/Y _5093_/X _5109_/X _5110_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_3_880 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_891 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_907 VGND VPWR sky130_fd_sc_hd__decap_8
X_5041_ _5036_/Y _5040_/X _5041_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_100_918 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4495__A _4492_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_169 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2727__B _2728_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_802 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_898 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_228 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3915__A2_N _3914_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_194 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_345 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_751 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_902 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3839__A _3839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2743__A _2719_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_929 VGND VPWR sky130_fd_sc_hd__decap_6
X_4825_ _4822_/X _4825_/B _4832_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5476__D _5476_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_4756_ _4756_/A _3778_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_3707_ _3727_/A _3687_/X _3707_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4687_ _4674_/A _4687_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_135_826 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_111 VGND VPWR sky130_fd_sc_hd__decap_8
X_3638_ _5284_/Y _3638_/B _3666_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_49_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_133 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3293__B key_in[87] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_829 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_913 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4532__B1 mode VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_57 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_3569_ _3569_/A _3570_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3886__A2 _3864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5308_ _5264_/X _5307_/X _5270_/X _5308_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_130_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_756 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2918__A _2918_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5239_ _4817_/A _5238_/X _4817_/A _5238_/X _5239_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_117 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4835__A1 _4802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4835__B2 _4815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_589 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4599__B1 _4600_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4852__B _4851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_345 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_762 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_98 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3749__A _3739_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_367 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_913 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_212 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_890 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_234 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_907 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_245 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3810__A2 _3697_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_256 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_968 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_42 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_267 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5386__D _4771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_928 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5012__A1 _4996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5372__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_428 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_289 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_776 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_427 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4220__C1 _4219_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_962 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3574__A1 _5178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4771__B1 data_out1[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_837 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3484__A _3484_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2782__C1 _2781_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5315__A2 _5313_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_655 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_509 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_445 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5079__B2 _5078_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_850 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_916 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3931__B _3913_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2828__A _2828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4826__A1 _4802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_426 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4826__B2 _4815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5204__A _4618_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_459 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2837__B1 _2836_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_515 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_824 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5251__A1 data_in2[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_250 VGND VPWR sky130_fd_sc_hd__fill_2
X_2940_ _5497_/Q _3110_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_31_710 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_907 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2967__B1_N _2966_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2871_ _2871_/A _2871_/B _2871_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5264__B1_N _5241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5003__A1 _5000_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4610_ _4609_/X _4610_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_787 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_81 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_940 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3565__A1 _3564_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4541_ _4541_/A _4541_/B _4541_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4762__B1 data_out1[12] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3394__A _5537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_943 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_325 VGND VPWR sky130_fd_sc_hd__decap_8
X_4472_ _4475_/A _4472_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_7_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_155 VGND VPWR sky130_fd_sc_hd__fill_2
X_3423_ _3422_/X _3484_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4002__B _4001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3868__A2 _3867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_220 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_743 VGND VPWR sky130_fd_sc_hd__decap_4
X_3354_ _3354_/A _3309_/Y _3354_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4937__B _4928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_776 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_553 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_938 VGND VPWR sky130_fd_sc_hd__decap_8
X_3285_ _3170_/A _3285_/B _3285_/C _3285_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_97_286 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5114__A _4891_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_437 VGND VPWR sky130_fd_sc_hd__fill_2
X_5024_ _5562_/Q _5014_/X _5024_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_66_662 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_898 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_120 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_879 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5460__RESET_B _4410_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5242__A1 _5239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5395__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3569__A _3569_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3869__A2_N _3868_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3288__B _3285_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_4808_ _5448_/Q _4811_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_10_938 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4753__B1 data_out1[8] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2920__B _2920_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4739_ _5542_/Q _4736_/X data_out2[31] _4737_/X _4739_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_147_472 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_419 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_314 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_133 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_144 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3308__B2 _3318_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__B _5006_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3859__A2 _5530_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_426 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5024__A _5562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5548__RESET_B _4305_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_504 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4863__A _4863_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_470 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3492__B1 _3462_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_835 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_559 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_194 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_805 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3479__A _3478_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_507 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5233__B2 _5258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2814__C _2813_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3795__A1 _3773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3198__B _3196_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_40 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3547__A1 _3521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_450 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3926__B _3924_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4744__B1 data_out1[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_62 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_781 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4103__A _4077_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_678 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5313__A2_N _5322_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_452 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_518 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_829 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_881 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_497 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3942__A _3941_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_448 VGND VPWR sky130_fd_sc_hd__fill_2
X_3070_ _3069_/A _3068_/Y _3071_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_76_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_429 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3483__B1 _3540_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3389__A _3317_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_698 VGND VPWR sky130_fd_sc_hd__decap_4
X_3972_ _3972_/A _3971_/X _3972_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_51_849 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_704 VGND VPWR sky130_fd_sc_hd__fill_2
X_2923_ _2849_/A _2921_/X _2923_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4599__A2_N _4600_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_2854_ _2733_/A _2698_/B _2876_/A _2854_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_164_707 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_269 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3538__B2 _3537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4735__B1 data_out2[29] VGND VPWR sky130_fd_sc_hd__diode_2
X_2785_ _2762_/Y _2770_/Y _2761_/Y _2785_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_5573_ _4573_/X _4573_/A _4274_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_163_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5109__A _5082_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_111 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_954 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4013__A _3180_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4524_ _4524_/A _4524_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_144_442 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_924 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_689 VGND VPWR sky130_fd_sc_hd__decap_12
X_4455_ _4469_/A _4461_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_177 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_136 VGND VPWR sky130_fd_sc_hd__fill_2
X_3406_ _3337_/A key_in[90] _3406_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4386_ _4387_/A _4386_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_905 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_916 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3171__C1 _3170_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3337_ _3337_/A key_in[88] _3337_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_501 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_735 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_234 VGND VPWR sky130_fd_sc_hd__decap_8
X_3268_ _5469_/Q _3266_/B _3267_/Y _3268_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_58_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_578 VGND VPWR sky130_fd_sc_hd__fill_2
X_5007_ _5008_/A _5006_/Y _5007_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3474__B1 _3472_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3199_ _3199_/A _3198_/Y _3199_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_26_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_194 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2915__B _2914_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_131 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5215__B2 _5226_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_484 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3777__B2 _3776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_534 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2931__A _2905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_99 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3746__B _3744_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_943 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5019__A _5002_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5410__CLK _5402_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_65 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_784 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_934 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3762__A _3749_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2_0_clock_A clkbuf_2_3_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_76 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5151__B1 _5143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4577__B _4576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_478 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_562 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_873 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5560__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5382__RESET_B _4502_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_779 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4257__A2 _4667_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_150 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_738 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_835 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_481 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_194 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_334 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2825__B key_in[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3002__A _2790_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3359__D _3358_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_871 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3937__A _3937_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_595 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_729 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4717__B1 data_out2[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_781 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5574__D _4574_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_954 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4193__B2 _4192_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_751 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4948__B1_N _4947_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_773 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3940__A1 _3939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_998 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_794 VGND VPWR sky130_fd_sc_hd__decap_3
X_4240_ _4222_/X _4227_/X _3848_/X _4244_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__5142__B1 _5128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1011 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_670 VGND VPWR sky130_fd_sc_hd__decap_12
X_4171_ _4073_/X _4170_/X _4171_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_68_746 VGND VPWR sky130_fd_sc_hd__fill_1
X_3122_ _4638_/X _3118_/X _3119_/X _3120_/X _3121_/X _3122_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_110_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_705 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4248__A2 _3788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_587 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_738 VGND VPWR sky130_fd_sc_hd__fill_2
X_3053_ _2973_/Y _3006_/X _3052_/X _3057_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_82_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_790 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_602 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3512__B1_N _3540_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_462 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_473 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_624 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4008__A _3983_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3955_ _5534_/Q _3955_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4950__B _4949_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_167 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_534 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_189 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2751__A _2750_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2906_ _4642_/A _2903_/B _2905_/Y _2913_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3527__B1_N _3526_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3886_ _3861_/X _3864_/Y _3860_/X _3886_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__5433__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4708__B1 data_out2[15] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_504 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2982__A2 _2981_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2837_ _2770_/Y _2834_/X _2836_/Y _2837_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__5484__D _3677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4184__A1 data_in1[27] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3285__C _3285_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_5556_ _4553_/X _4553_/A _4295_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2768_ _5334_/X _2769_/A _2767_/Y _2768_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_133_902 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_913 VGND VPWR sky130_fd_sc_hd__fill_2
X_4507_ _4504_/X _4507_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_272 VGND VPWR sky130_fd_sc_hd__decap_3
X_5487_ _3747_/X _5261_/A _4378_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2699_ _2885_/A _2852_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3582__A _4537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_434 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5133__B1 _5132_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4438_ _4438_/A _4438_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_618 VGND VPWR sky130_fd_sc_hd__fill_1
X_4369_ _4397_/A _4375_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4892__C1 _4891_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5005__C _4980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_407 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2926__A _2925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3447__B1 _3445_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_237 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5302__A _5301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_963 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_974 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_10 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_760 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5021__B _5019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_698 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_484 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_43 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_495 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_988 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_156 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_98 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_871 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_707 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_31 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_375 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_910 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5394__D _4787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4175__A1 _4172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1000 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2725__A2 _2691_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4588__A _3465_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5563__RESET_B _4287_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_307 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3686__B1 _3663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_36 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3150__A2 _3146_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_256 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_6_0_clock_A clkbuf_3_6_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_418 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_598 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3623__A2_N _3622_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_749 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3989__A1 _3939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_142 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5569__D _5569_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_451 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_771 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_782 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_635 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5456__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3667__A _3666_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_487 VGND VPWR sky130_fd_sc_hd__fill_2
X_3740_ _5292_/X _3738_/X _3739_/Y _3740_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_159_887 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_718 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_515 VGND VPWR sky130_fd_sc_hd__decap_4
X_3671_ _3671_/A _3670_/X _3671_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5191__A2_N _5190_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_537 VGND VPWR sky130_fd_sc_hd__decap_8
X_5410_ _5410_/D data_out2[8] _4470_/X _5402_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4166__A1 data_in1[26] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5363__B1 _5331_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_913 VGND VPWR sky130_fd_sc_hd__fill_2
X_5341_ _4848_/A _5341_/B _2769_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_127_784 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4498__A _4501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_732 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5115__B1 _4942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_808 VGND VPWR sky130_fd_sc_hd__decap_12
X_5272_ _5264_/X _5271_/X _5264_/X _5271_/X _5272_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_141_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_4223_ _3395_/X _3521_/X _3395_/X _3521_/X _4225_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3677__B1 _3654_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_4154_ _4151_/X _4153_/Y _4151_/X _4153_/Y _4154_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_565 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4945__B _4944_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3105_ _5529_/Q _3133_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4085_ _4784_/X _4083_/X _4115_/B _4113_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__2746__A _2745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5122__A _5122_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3451__B1_N _3450_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3036_ _2966_/A _3036_/B _2965_/Y _3036_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_36_451 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5479__D _3580_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4641__A2 _4631_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_613 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4961__A _4961_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_495 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_646 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_117 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_465 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_128 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4987_ _4987_/A _4986_/X _4987_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_11_318 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__A _3577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_331 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3938_ _3931_/X _3937_/X _3938_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_137_504 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3296__B _3295_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2955__A2 _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_846 VGND VPWR sky130_fd_sc_hd__fill_2
X_3869_ _3866_/X _3868_/Y _3866_/X _3868_/Y _3869_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5354__B1 _5321_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_740 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_5539_ _5539_/D _5539_/Q _4315_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_423 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3380__A2 _3379_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4201__A _4195_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_968 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_927 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_798 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_949 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_521 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_830 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_841 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4855__B _4854_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_930 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_749 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5032__A _5031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_183 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_941 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5479__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_194 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_440 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_451 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5389__D _4776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_64 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4871__A _4871_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_605 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A3 _5184_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__A _3426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_796 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_830 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_504 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_13_0_clock_A clkbuf_3_6_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_85 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4148__A1 _4100_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4148__B2 _4131_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_740 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_867 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_355 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_762 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_209 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_890 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_592 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5207__A _5207_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_540 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3371__A2 _3369_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3659__B1 _3588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3950__A _3839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_800 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_971 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2882__A1 data_in2[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_387 VGND VPWR sky130_fd_sc_hd__decap_8
X_4910_ _5553_/Q _4909_/X _5553_/Q _4909_/X _4910_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4781__A _4672_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_292 VGND VPWR sky130_fd_sc_hd__decap_4
X_4841_ _4840_/A _4839_/X _4840_/X _4841_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3397__A _5510_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_4772_ _2889_/A _3113_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_802 VGND VPWR sky130_fd_sc_hd__decap_3
X_3723_ _2735_/X _3722_/X _3723_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_146_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4005__B _3984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4139__A1 _4788_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3654_ _3615_/A _3570_/B _5327_/A _3654_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5485__RESET_B _4380_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_378 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3844__B _3843_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_721 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5414__RESET_B _4465_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3585_ _3585_/A _3586_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_127_592 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5117__A _5569_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_5324_ _5256_/A _5323_/X _5324_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__4021__A _4016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_905 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_509 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_616 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2771__A2_N _2770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_798 VGND VPWR sky130_fd_sc_hd__fill_2
X_5255_ _5227_/B _5254_/Y _5256_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_735 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4956__A _4921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3860__A _3750_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_852 VGND VPWR sky130_fd_sc_hd__fill_2
X_4206_ _4187_/B _4192_/Y _4073_/X _4212_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3114__A2 _3088_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_800 VGND VPWR sky130_fd_sc_hd__decap_8
X_5186_ _4635_/A _5207_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_68_373 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_4137_ _4130_/X _4136_/Y _4130_/X _4136_/Y _4137_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_226 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2873__B2 _2872_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4068_ _4068_/A _4066_/X _4069_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_56_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_782 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_229 VGND VPWR sky130_fd_sc_hd__decap_3
X_3019_ _3020_/A _3020_/B _3021_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_24_410 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_977 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2923__B _2921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_605 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_115 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_947 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3100__A _2927_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2928__A2 _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_159 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_172 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_857 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_55 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_304 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_378 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3754__B _3734_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_37 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_859 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5027__A _5027_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_702 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_381 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4866__A _4852_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_54 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3770__A _4707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_800 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_256 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_971 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_982 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4853__A2 _4851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_237 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_74 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_814 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4066__B1 _4065_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_549 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_977 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3929__B _3812_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_402 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_785 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_498 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__A _4102_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_971 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3010__A _3010_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_982 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2919__A2 _2918_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_621 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3945__A _3945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_120 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_697 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4245__A2_N _4244_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3370_ _3178_/Y _3369_/X _3370_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_713 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_81 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_947 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_735 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_392 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_446 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3680__A _3680_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5040_ _5564_/Q _5039_/X _5564_/Q _5039_/X _5040_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_790 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4057__B1 _3273_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_207 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_387 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3839__B _3812_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_368 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_914 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_251 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2743__B _2718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_571 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_908 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_947 VGND VPWR sky130_fd_sc_hd__decap_8
X_4824_ _4822_/X _4825_/B _4824_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__4016__A _3968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_301 VGND VPWR sky130_fd_sc_hd__decap_4
X_4755_ _3759_/A _4745_/X data_out1[9] _4746_/X _4755_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_147_643 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3855__A _3835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_654 VGND VPWR sky130_fd_sc_hd__fill_2
X_3706_ _3704_/X _3705_/Y _3706_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4686_ _5517_/Q _5356_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3454__A2_N _3464_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_186 VGND VPWR sky130_fd_sc_hd__fill_2
X_3637_ _5178_/Y _5520_/Q _3573_/A _3636_/Y _3638_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__5492__D _5492_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_903 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4532__B2 _4531_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3568_ _4664_/X _3569_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_1_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_702 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_69 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_925 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_936 VGND VPWR sky130_fd_sc_hd__fill_2
X_5307_ _4827_/A _5270_/B _5307_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_510 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4686__A _5517_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_690 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_3499_ _3499_/A _3528_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_5238_ _4636_/A _5234_/X _5235_/X _5236_/X _5237_/X _5238_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_130_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_660 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2918__B _2918_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4835__A2 _4842_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_68 VGND VPWR sky130_fd_sc_hd__decap_8
X_5169_ _5169_/A _5169_/B _5170_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_56_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_803 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4048__B1 _5529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_836 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_173 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2934__A _2934_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4599__B2 _4600_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5310__A _5309_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_357 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3749__B _3744_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_202 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5517__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_10 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_919 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_246 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_284 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_593 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_257 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_54 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5012__A2 _4995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_279 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4220__B1 _4205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_941 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3765__A _3765_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_991 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3574__A2 _3572_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4771__A1 _3902_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4771__B2 _4770_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2782__B1 _2733_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3484__B _3457_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_635 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_634 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3594__A1_N _3583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_166 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4596__A _4595_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_690 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3297__B1_N _3296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_40 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_862 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_800 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4826__A2 _4824_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5204__B key_in[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_310 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_438 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2837__A1 _2770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_641 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3005__A _3004_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_527 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2844__A _2855_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5251__A2 _5222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_677 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5577__D _4260_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_295 VGND VPWR sky130_fd_sc_hd__fill_2
X_2870_ _2870_/A _2870_/B _2871_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_31_755 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5003__A2 _4999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4211__B1 _3508_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_287 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3675__A _3674_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4540_ _4837_/B _4541_/B _4540_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_129_665 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4762__A1 _2714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3565__A2 _3564_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_900 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4762__B2 _4758_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_816 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_984 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_304 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2773__B1 _2736_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4471_ _4475_/A _4471_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_128_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_955 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_337 VGND VPWR sky130_fd_sc_hd__decap_3
X_3422_ _3395_/X _3421_/X _3422_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_171_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_3353_ _3353_/A _3356_/B _3359_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_98_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_405 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_928 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_565 VGND VPWR sky130_fd_sc_hd__decap_12
X_3284_ _3284_/A _3282_/X _3285_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_57_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5114__B _5114_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5023_ _5023_/A _5027_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_298 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_855 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_877 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_888 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_674 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_460 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3818__B1_N _3817_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2754__A _5300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5130__A _5052_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_132 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5242__A2 _5241_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3789__C1 _3788_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5487__D _3747_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_688 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4137__A2_N _4136_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5053__A1_N _5065_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_593 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_48 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_744 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_4807_ _4798_/X _4813_/A _4802_/X _4798_/B _4806_/X _4807_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_166_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_941 VGND VPWR sky130_fd_sc_hd__decap_4
X_2999_ _2999_/A _2999_/B _2999_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3585__A _3585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4753__A1 _5261_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4738_ _5541_/Q _4736_/X data_out2[30] _4737_/X _5432_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4753__B2 _4746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_421 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_955 VGND VPWR sky130_fd_sc_hd__decap_4
X_4669_ _4631_/Y _4662_/Y _3676_/A _4668_/Y _4669_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_163_977 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_510 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2929__A _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_34 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_744 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_659 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_874 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_576 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_587 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5024__B _5014_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_65 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4863__B _4862_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_516 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3492__A1 data_in2[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_700 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5397__D _4792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5517__RESET_B _4342_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2814__D _2814_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3198__C _3197_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3795__A2 _3774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_563 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3495__A _3178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_247 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4744__A1 _5260_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3547__A2 _3537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4744__B2 _4737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_270 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_860 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_638 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_497 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_825 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3483__A1 _3463_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4680__B1 data_out2[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_836 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_655 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_677 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3389__B _3389_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_3971_ _3968_/X _3970_/Y _3971_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_44_880 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_198 VGND VPWR sky130_fd_sc_hd__decap_12
X_2922_ _2849_/B _2921_/X _2924_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_93_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_2853_ data_in2[10] _2731_/X _2812_/X _2852_/Y _2853_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_31_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_440 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4735__A1 _3493_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_5572_ _4572_/X _4572_/A _4277_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4735__B2 _4726_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2784_ _2784_/A _2779_/Y _2784_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_117_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_782 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5109__B _5109_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4523_ _4523_/A _4578_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4013__B _4012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_977 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_145 VGND VPWR sky130_fd_sc_hd__decap_8
X_4454_ _4449_/A _4454_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_936 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_947 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3742__B1_N _3741_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3405_ _3337_/A key_in[26] _3405_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2749__A _2718_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_969 VGND VPWR sky130_fd_sc_hd__decap_12
X_4385_ _4387_/A _4385_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_852 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3171__B1 _3143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5125__A _5125_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_563 VGND VPWR sky130_fd_sc_hd__decap_4
X_3336_ _3293_/A key_in[24] _3336_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_58_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_928 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_874 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_939 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_747 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4964__A _5462_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3267_ _3344_/A _3267_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3439__A1_N _4784_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5006_ _4988_/X _5004_/X _5005_/X _5006_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_27_814 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3474__A1 _4640_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_162 VGND VPWR sky130_fd_sc_hd__fill_2
X_3198_ _3195_/X _3196_/X _3197_/Y _3198_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_66_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3474__B2 _3473_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_324 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_655 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_666 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_891 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_894 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2931__B _2913_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_760 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3746__C _3745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_729 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5019__B _5019_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_635 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2951__B1_N _2950_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_251 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_679 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_167 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_638 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3762__B _3782_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5151__A1 _4857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5151__B2 _4815_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_957 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_979 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3162__B1 _3154_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_21 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_416 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_395 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_54 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4874__A _4874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_205 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_869 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_806 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_305 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_828 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_880 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3002__B key_in[79] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_390 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_541 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_51 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3937__B _3936_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4717__A1 _3175_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4114__A _4065_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4717__B2 _4713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_578 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_966 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3953__A _3939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_977 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3940__A2 _3904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_487 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_638 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5142__A1 _4857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5385__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5142__B2 _4815_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4154__A1_N _4151_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3238__A2_N _3237_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3153__B1 _3124_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_4170_ _4152_/A _4136_/Y _4093_/X _4170_/D _4170_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_110_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_991 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_682 VGND VPWR sky130_fd_sc_hd__decap_3
X_3121_ _3043_/X key_in[114] _3044_/X _3121_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_95_533 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4784__A _3108_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_866 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4248__A3 _5510_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_3052_ _3052_/A _3052_/B _3052_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_899 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5439__RESET_B _4435_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_633 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_817 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_839 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_794 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4008__B _4008_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_891 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_3954_ _3904_/X _3953_/X _3954_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_502 VGND VPWR sky130_fd_sc_hd__decap_12
X_2905_ _2905_/A _2905_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_31_371 VGND VPWR sky130_fd_sc_hd__fill_2
X_3885_ _3794_/A _3884_/X _3885_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__4708__A1 _3020_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_579 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4708__B2 _4701_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2836_ _2761_/A _2835_/X _2794_/X _2836_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__4024__A _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_549 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4184__A2 _4125_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5555_ _4552_/X _4944_/A _4296_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2767_ _2767_/A _2767_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3863__A _3818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_977 VGND VPWR sky130_fd_sc_hd__fill_1
X_4506_ _4504_/X _4506_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_925 VGND VPWR sky130_fd_sc_hd__decap_12
X_5486_ _3718_/X _5229_/A _4379_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2698_ _5252_/A _2698_/B _5518_/Q _2698_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5133__A1 _5132_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4437_ _4438_/A _4437_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_132_446 VGND VPWR sky130_fd_sc_hd__decap_12
X_4368_ _4367_/A _4368_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4892__B1 _4531_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_533 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4694__A _5521_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3319_ _3465_/A _3319_/B _3320_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_101_855 VGND VPWR sky130_fd_sc_hd__decap_8
X_4299_ _4303_/A _4299_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_877 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3447__A1 _4640_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_739 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2926__B _2924_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_611 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3447__B2 _3446_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_920 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5302__B key_in[68] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_644 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_79 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_655 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3103__A _3026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_817 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_22 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5312__A2_N _5311_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_33 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_349 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_66 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_800 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2942__A _2943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_833 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_321 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_883 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_343 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_382 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_719 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_544 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_43 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_54 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_229 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4175__A2 _4174_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_977 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3383__B1 _3373_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4588__B _4588_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1004 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_413 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_733 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3686__A1 _3661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_371 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4883__B1 _4873_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_235 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3150__A3 _3147_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_706 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_268 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_503 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5532__RESET_B _4324_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3989__A2 _3988_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_655 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_964 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_750 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3013__A _3012_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_50 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2852__A _2852_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2949__B1 _2998_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_855 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3610__A1 _3583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_382 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3162__A2_N _3161_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_899 VGND VPWR sky130_fd_sc_hd__decap_12
X_3670_ _3658_/Y _3669_/X _3670_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_9_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_549 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4166__A2 _4125_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5363__A1 _5325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_903 VGND VPWR sky130_fd_sc_hd__decap_4
X_5340_ _4636_/A _5336_/X _5337_/X _5338_/X _5339_/X _5341_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_56_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_593 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5115__A1 _5473_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_5271_ _4827_/A _5270_/B _5270_/X _5271_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_114_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_4222_ _3848_/X _4211_/X _4212_/A _4222_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_99_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_265 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3677__A1 data_in1[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_820 VGND VPWR sky130_fd_sc_hd__decap_4
X_4153_ _4073_/X _4152_/X _4095_/X _4153_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_68_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_352 VGND VPWR sky130_fd_sc_hd__fill_2
X_3104_ _2885_/A _3170_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_205 VGND VPWR sky130_fd_sc_hd__decap_12
X_4084_ _4784_/X _4083_/X _4115_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5122__B _5138_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_953 VGND VPWR sky130_fd_sc_hd__fill_2
X_3035_ _3015_/A _3014_/A _3037_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_36_430 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4019__A _3970_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5400__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_463 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_772 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_219 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4961__B _4960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_945 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3858__A _5530_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_433 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_619 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_4986_ _4997_/C _4976_/X _4975_/X _4986_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__B _3600_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3937_ _3937_/A _3936_/X _3937_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XANTENNA__5495__D _3928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5550__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_814 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_516 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_302 VGND VPWR sky130_fd_sc_hd__fill_2
X_3868_ _3794_/A _3867_/X _3815_/Y _3868_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_20_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5354__A1 data_in2[5] VGND VPWR sky130_fd_sc_hd__diode_2
X_2819_ _2819_/A _2819_/B _2872_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_3799_ _3797_/X _3799_/B _3799_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_560 VGND VPWR sky130_fd_sc_hd__fill_2
X_5538_ _5538_/D _5538_/Q _4316_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_947 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4201__B _4232_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_5469_ _5063_/X _5469_/Q _4399_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_552 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_766 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_39 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_276 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4865__B1 _4864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_691 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_34 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_641 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2937__A _4943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_419 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3240__A1_N _3249_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_385 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_696 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_290 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_260 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_794 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_422 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__A _3681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_764 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__B _3485_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_179 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_140 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_190 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_685 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_516 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_858 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_846 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4148__A2 _4132_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_879 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_345 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_574 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_788 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3823__A1_N _2914_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_596 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3659__B2 _5521_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3950__B _3950_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2847__A _2847_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_330 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_490 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_341 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5223__A _5223_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5423__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2882__A2 _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4608__B1 _4607_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_249 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_400 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_934 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5573__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3678__A _4664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_731 VGND VPWR sky130_fd_sc_hd__fill_1
X_4840_ _4840_/A _4839_/X _4840_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_61_786 VGND VPWR sky130_fd_sc_hd__decap_3
X_4771_ _3902_/C _4769_/X data_out1[16] _4770_/X _4771_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3722_ _5284_/Y _5524_/Q _5515_/Q _3721_/Y _3722_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_159_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_195 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4139__A2 _4137_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3653_ data_in1[4] _3581_/X _3633_/X _3652_/X _3653_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_162_806 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_357 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3347__B1 _3342_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4302__A _4303_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3584_ _4524_/Y _3584_/B _3585_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_5323_ _5285_/X _5322_/Y _5323_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5117__B _5101_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_541 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4021__B _4020_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_552 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_766 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_5254_ _5243_/X _5254_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_87_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4956__B _4955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5454__RESET_B _4417_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3860__B _3859_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4205_ _4126_/X _4090_/X _4794_/X _4205_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_5185_ _4618_/A key_in[64] _5185_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_812 VGND VPWR sky130_fd_sc_hd__decap_4
X_4136_ _3382_/X _4135_/X _3382_/X _4135_/X _4136_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_110_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_238 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_856 VGND VPWR sky130_fd_sc_hd__decap_8
X_4067_ _4068_/A _4066_/X _4069_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4972__A _4971_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5272__B1 _5264_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3018_ _2999_/Y _3017_/X _2999_/Y _3017_/X _3020_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_731 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3588__A _3588_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_1003 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4969_ _3052_/A _4968_/B _4968_/X _4971_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3100__B _3098_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_814 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_644 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_154 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3338__B1 _3222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4212__A _4212_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_327 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_49 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5027__B _5027_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_359 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5446__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_585 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4866__B _4855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_66 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5043__A _5036_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_823 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_21 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_493 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_867 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4882__A _4882_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4066__A1 _4021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_506 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5263__B1 _5262_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_377 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_411 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_720 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3194__A1_N _5023_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_591 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3929__C _3113_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_572 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_96 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__B _4105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_471 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_650 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_110 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3945__B _3945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_346 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_665 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5218__A _5192_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4122__A _4112_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_676 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3132__A1_N _3107_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_861 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_703 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_585 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4829__B1 _4542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_747 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3680__B _3669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3777__A1_N _3768_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_780 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_750 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4057__B2 _4056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_697 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_794 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_399 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_731 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3839__C _3875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_926 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_4823_ _4823_/A _4823_/B _4825_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_22_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_274 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3403__B1_N _3402_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4016__B _4019_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_611 VGND VPWR sky130_fd_sc_hd__fill_2
X_4754_ _5288_/A _3759_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_159_482 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_622 VGND VPWR sky130_fd_sc_hd__fill_2
X_3705_ _2723_/A _3703_/X _3705_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_30_992 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3855__B _3853_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4685_ _5321_/C _4674_/X data_out2[5] _4677_/X _5407_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_135_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5128__A _5128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_3636_ _5520_/Q _3636_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_134_316 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5469__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4032__A _4002_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_809 VGND VPWR sky130_fd_sc_hd__decap_12
X_3567_ _3564_/X _3565_/Y _3566_/Y _3567_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_115_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_872 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3871__A _3870_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5306_ _4836_/A _5334_/B _4836_/A _5334_/B _5306_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__3740__B1 _3739_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_371 VGND VPWR sky130_fd_sc_hd__fill_2
X_3498_ _3496_/X _3497_/X _3496_/X _3497_/X _3498_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_544 VGND VPWR sky130_fd_sc_hd__decap_6
X_5237_ _5234_/A key_in[98] _5303_/A _5237_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_102_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_503 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4835__A3 _4834_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5168_ _5169_/A _5169_/B _5170_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_96_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_642 VGND VPWR sky130_fd_sc_hd__decap_4
X_4119_ _4020_/Y _4119_/B _4119_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_57_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_664 VGND VPWR sky130_fd_sc_hd__decap_12
X_5099_ _4896_/X _5097_/X _5098_/Y _5090_/Y _4806_/X _5099_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XANTENNA__4048__A1 _3133_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4048__B2 _4047_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_325 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2934__B key_in[77] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_230 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4207__A _4000_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_550 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_203 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_775 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_786 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_225 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_274 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_959 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_258 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3559__B1 _3526_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_407 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2950__A _2989_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_622 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4220__A1 data_in1[29] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_99 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3765__B _3679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_441 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4771__A2 _4769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2939__A1_N _2931_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_975 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_452 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_603 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5038__A _5563_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2782__A1 data_in2[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_165 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_176 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_647 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5376__RESET_B _4509_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4877__A _4875_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_861 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_552 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_679 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_403 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3731__B1 _3730_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_52 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_812 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4826__A3 _4832_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2837__A2 _2834_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_667 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_230 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4117__A _4063_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3021__A _3021_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_881 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_745 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4133__B1_N _4132_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2860__A _2861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_255 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_72 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_791 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4211__B2 _4210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__B _3674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_964 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4762__A2 _4757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_440 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_912 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2773__B2 _2772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3970__B1 _3969_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4470_ _4475_/A _4470_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_316 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_198 VGND VPWR sky130_fd_sc_hd__decap_12
X_3421_ _3436_/A _3420_/Y _3436_/A _3420_/Y _3421_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3722__B1 _5515_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_511 VGND VPWR sky130_fd_sc_hd__decap_8
X_3352_ _3284_/A _3352_/B _3356_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_124_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_853 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_190 VGND VPWR sky130_fd_sc_hd__fill_2
X_3283_ _3284_/A _3282_/X _3285_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_140_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_577 VGND VPWR sky130_fd_sc_hd__decap_3
X_5022_ _4896_/X _5020_/X _5021_/Y _5017_/A _4806_/X _5022_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_85_428 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5114__C _5114_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_804 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_837 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_196 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2754__B key_in[40] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5130__B _5130_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3789__B1 _3765_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_667 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4027__A _4013_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_200 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_717 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2770__A _2770_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_918 VGND VPWR sky130_fd_sc_hd__fill_2
X_4806_ _4815_/A _4806_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2998_ _2998_/A _2998_/B _2998_/C _2887_/X _2999_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_9_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4753__A2 _4745_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4737_ _4701_/A _4737_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_452 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3669__A1_N _3665_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_625 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3961__B1 _3960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_102 VGND VPWR sky130_fd_sc_hd__decap_12
X_4668_ _4667_/X _4668_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_162_433 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_198 VGND VPWR sky130_fd_sc_hd__fill_2
X_3619_ _3619_/A _3619_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4599_ _4600_/A _4600_/B _4600_/A _4600_/B _4599_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_162_477 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_308 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_211 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2929__B _2884_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_244 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_28 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_599 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_620 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_439 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_322 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_962 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3607__A1_N _3601_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2945__A _2945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_815 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5321__A _5252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_601 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3492__A2 _3391_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_612 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_848 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_678 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_745 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_216 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_586 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5557__RESET_B _4294_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3495__B _3495_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4744__A2 _4736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_259 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_282 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_988 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_91 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4400__A _4402_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_211 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_428 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2855__A _2855_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_83 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5209__B1 _5205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_910 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4680__A1 _4679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_995 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3483__A2 _3482_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4680__B2 _4677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3453__A2_N _3452_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_848 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_100 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2691__B1 _5358_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3389__C _3388_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_3970_ _3918_/Y _3943_/X _3969_/X _3970_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_50_317 VGND VPWR sky130_fd_sc_hd__fill_2
X_2921_ _2850_/A _2921_/B _2921_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_728 VGND VPWR sky130_fd_sc_hd__decap_4
X_2852_ _2852_/A _2855_/B _2851_/X _2852_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_148_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_586 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_249 VGND VPWR sky130_fd_sc_hd__fill_2
X_5571_ _4571_/X _5571_/Q _4278_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2783_ _2733_/A _2698_/B _2847_/A _2783_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_129_452 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4735__A2 _4725_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_4522_ _4522_/A _4523_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_157_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_422 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1007 VGND VPWR sky130_fd_sc_hd__decap_12
X_4453_ _4449_/A _4453_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3404_ _3334_/X key_in[58] _3404_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4010__B1_N _4009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4310__A _4305_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4384_ _4387_/A _4384_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_520 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2749__B _2743_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3171__A1 data_in2[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_149 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5125__B _5124_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3335_ _3334_/X key_in[56] _3335_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5507__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_214 VGND VPWR sky130_fd_sc_hd__fill_2
X_3266_ _5469_/Q _3266_/B _3344_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_86_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_5005_ _4982_/A _4992_/A _4980_/X _5005_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__2765__A _5345_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3197_ _3125_/Y _3197_/B _3129_/Y _3197_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__5141__A _5148_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3474__A2 _3470_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_921 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_483 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5498__D _5498_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4967__A1_N _4555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4980__A _4968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3593__A1_N _3587_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_520 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_24 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3596__A _3596_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_748 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_923 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_978 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_466 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5316__A _5276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_105 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_499 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5151__A2 _5149_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_413 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_680 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_947 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3162__B2 _3161_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1018 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_886 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_737 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_439 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4874__B _4873_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4111__B1 _4095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_450 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5051__A _5564_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_770 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_280 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_645 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_965 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_144 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4890__A _4886_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_818 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_513 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5391__RESET_B _4492_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4717__A2 _4712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_901 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4114__B _4117_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_422 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_433 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3953__B _3952_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_989 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_763 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_797 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5226__A _5226_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_785 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_436 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5142__A2 _5139_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_458 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3153__A1 _3125_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_190 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4136__A2_N _4135_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_812 VGND VPWR sky130_fd_sc_hd__decap_12
X_3120_ _3077_/A key_in[82] _3120_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_160 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_490 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_962 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4102__B1 _4101_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_409 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_3051_ _2977_/Y _3050_/X _3051_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_83_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_601 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_770 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_239 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5067__A1_N _5566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_494 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_987 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_261 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4008__C _4006_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5479__RESET_B _4387_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1011 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_125 VGND VPWR sky130_fd_sc_hd__decap_12
X_3953_ _3939_/X _3952_/X _3953_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_50_147 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5408__RESET_B _4472_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_514 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2967__A1 _2966_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4305__A _4305_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2904_ _2904_/A _2905_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_3884_ _3823_/X _3847_/X _3866_/X _3814_/X _3884_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_149_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_558 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4708__A2 _4699_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2835_ _4900_/A _2794_/B _2835_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_394 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4024__B _4027_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_923 VGND VPWR sky130_fd_sc_hd__decap_8
X_2766_ _2766_/A _2767_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_5554_ _5554_/D _5554_/Q _4298_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3863__B _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4505_ _4504_/X _4505_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_455 VGND VPWR sky130_fd_sc_hd__fill_2
X_5485_ _3696_/X _5200_/A _4380_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2697_ data_in2[6] _5222_/X _5356_/X _2696_/X _5517_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_144_252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_937 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5136__A _5110_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_583 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4040__A _4039_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_4436_ _4438_/A _4436_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5133__A2 _5131_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_4367_ _4367_/A _4367_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4975__A _4921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_361 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4892__A1 _4882_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_672 VGND VPWR sky130_fd_sc_hd__fill_2
X_3318_ _3318_/A _3318_/B _3319_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_101_834 VGND VPWR sky130_fd_sc_hd__fill_2
X_4298_ _4303_/A _4298_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_867 VGND VPWR sky130_fd_sc_hd__decap_4
X_3249_ _3248_/Y _3249_/B _3176_/X _3249_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_67_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_589 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_36 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3447__A2 _3443_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_111 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_740 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3103__B _3143_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_667 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_998 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_34 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_45 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_659 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2942__B _2943_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_979 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_812 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4215__A _4214_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3080__B1 _3078_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_895 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_394 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_208 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_33 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_539 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_527 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_422 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_509 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_904 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3383__B2 _3382_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4229__A1_N _3523_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5046__A _5047_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1016 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_285 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_458 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4885__A _4885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_288 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4883__A1 _4874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3686__A2 _3667_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_299 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_225 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_81 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3188__B1_N _3187_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_634 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_943 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3013__B _3012_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_762 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_166 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3111__B1_N _3160_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5572__RESET_B _4277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_648 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2852__B _2855_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5501__RESET_B _4360_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_834 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2949__B2 _2948_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4125__A _4533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_361 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3610__A2 _3593_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5363__A2 _5332_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_572 VGND VPWR sky130_fd_sc_hd__decap_8
X_5270_ _4827_/A _5270_/B _5270_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5115__A2 _4995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_593 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VPWR sky130_fd_sc_hd__decap_8
X_4221_ _4126_/X _3569_/A _3368_/A _4221_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_123_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_277 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3677__A2 _3581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_299 VGND VPWR sky130_fd_sc_hd__fill_2
X_4152_ _4152_/A _4136_/Y _4152_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_854 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_556 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_3103_ _3026_/A _3143_/B _5529_/Q _3103_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_56_707 VGND VPWR sky130_fd_sc_hd__fill_1
X_4083_ _4075_/Y _4082_/X _4075_/Y _4082_/X _4083_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_898 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_397 VGND VPWR sky130_fd_sc_hd__fill_2
X_3034_ _3032_/A _3032_/B _3033_/Y _3038_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4019__B _4019_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_965 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_209 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_968 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4643__A2_N _4641_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_4985_ _5464_/Q _4985_/X VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3936_ _3075_/Y _3933_/X _3935_/X _3936_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_51_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_990 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_3867_ _3823_/X _3847_/X _3867_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_137_528 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3874__A _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_325 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_859 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5354__A2 _5222_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2818_ _5361_/A _3895_/A _4750_/X _3012_/A _2819_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_3798_ _3682_/Y _3796_/X _3799_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_164_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_36 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_764 VGND VPWR sky130_fd_sc_hd__fill_2
X_5537_ _5537_/D _5537_/Q _4317_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2749_ _2718_/B _2743_/Y _2749_/C _2748_/Y _2749_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_145_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_200 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_520 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5277__B1_N _5276_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5468_ _5048_/Y _5468_/Q _4400_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3117__A1 _3116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_778 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_575 VGND VPWR sky130_fd_sc_hd__decap_4
X_4419_ _4419_/A _4422_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4865__A1 _4863_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5399_ _5399_/D data_out1[29] _4482_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_597 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3299__A2_N _3298_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_480 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2937__B _2936_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_559 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2953__A _2930_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_114 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_434 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3768__B _3767_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_108 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5375__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_158 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3237__A2_N _3236_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3053__B1 _3052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_43 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_21 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_821 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_990 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_32 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_675 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_152 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_803 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_174 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_314 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_876 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_825 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_313 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_196 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_375 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4148__A3 _4107_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_509 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_117 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_428 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3950__C _5497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2847__B _2847_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_824 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4608__A1 _4646_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3024__A _2927_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_921 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_879 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3959__A _3909_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_721 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_957 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_253 VGND VPWR sky130_fd_sc_hd__decap_12
X_4770_ _4700_/A _4770_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_3721_ _5524_/Q _3721_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4792__B1 data_out1[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_697 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_837 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3694__A _3694_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_3652_ _3579_/A _3650_/Y _3651_/X _3652_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_162_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3347__B2 _3346_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_3583_ _3615_/A _3570_/B _3583_/C _3583_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_161_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_881 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_5322_ _5322_/A _5322_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_6_891 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_778 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_873 VGND VPWR sky130_fd_sc_hd__decap_12
X_5253_ _5514_/Q _5253_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_102_428 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_832 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_4204_ data_in1[28] _4125_/X _4185_/X _4203_/Y _4204_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_5184_ _4618_/A key_in[0] _5184_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4135_ _4133_/X _4134_/X _4133_/X _4134_/X _4135_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_984 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_16 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5494__RESET_B _4370_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5326__A2_N _4756_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_4066_ _4021_/X _4063_/X _4065_/Y _4066_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_83_334 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4972__B _4970_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_49 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5398__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5423__RESET_B _4454_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5272__B2 _5271_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3017_ _3892_/A _3016_/X _3892_/A _3016_/X _3017_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_913 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3648__B1_N _3647_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_592 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1015 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_428 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_618 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4968_ _3052_/A _4968_/B _4968_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3100__C _3099_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4783__B1 data_out1[22] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3919_ _3032_/A _3917_/X _3918_/Y _3925_/A VGND VPWR sky130_fd_sc_hd__a21o_4
X_4899_ _5552_/Q _4899_/B _4899_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_137_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_818 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3338__A1 _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4212__B _4211_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_840 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_564 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_726 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5324__A _5256_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_748 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_640 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5043__B _5040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3161__A2_N _3160_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_995 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_194 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_879 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4066__A2 _4063_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5263__A1 _5260_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_762 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3779__A _3778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3274__B1 _3250_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_849 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_765 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_478 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_489 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_990 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_450 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_459 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4774__B1 data_out1[18] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_48 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_611 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4403__A _4402_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_684 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_358 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5218__B _5216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_550 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4122__B _4120_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_572 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3019__A _3020_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_188 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_125 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_61 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2858__A _2858_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5234__A _5234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4829__B2 _4828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_662 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5540__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_548 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_304 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_529 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3265__B1 _3263_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_337 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5006__A1 _4988_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4822_ _4821_/A _4821_/B _4821_/X _4822_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3017__B1 _3892_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_286 VGND VPWR sky130_fd_sc_hd__decap_12
X_4753_ _5261_/A _4745_/X data_out1[8] _4746_/X _4753_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_30_960 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_314 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4613__A1_N _5446_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3704_ _3603_/B _3703_/X _3704_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3855__C _3854_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4313__A _4312_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4684_ _5516_/Q _5321_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_818 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_829 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4032__B _4009_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3635_ _3586_/A _3634_/X _3635_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_146_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5190__B1 _5211_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3566_ _5197_/A _2852_/A _5542_/Q data_in2[31] _4546_/A _3566_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_89_916 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3740__A1 _5292_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5305_ _4637_/A _5300_/X _5301_/X _5302_/X _5304_/X _5334_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_142_361 VGND VPWR sky130_fd_sc_hd__decap_8
X_3497_ _3155_/Y _3466_/B _3466_/X _3468_/X _3497_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_737 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_5236_ _5236_/A key_in[66] _5236_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_124_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_651 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4983__A _4891_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5167_ _5167_/A _5167_/B _5169_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_68_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_537 VGND VPWR sky130_fd_sc_hd__fill_2
X_4118_ _4016_/X _4119_/B _4118_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_83_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_5098_ _5098_/A _5098_/B _5098_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_57_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4048__A2 _5538_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_367 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_816 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_676 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3599__A _3615_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4049_ _3932_/Y _4048_/X _4049_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_25_754 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4207__B _4097_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_204 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_242 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_916 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3008__B1 _2973_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_237 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3559__A1 _3396_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2950__B _2989_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_23 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_34 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_960 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4220__A2 _4125_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5319__A _5281_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_100 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_420 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_634 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3765__C _3778_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5413__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_492 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_987 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2782__A2 _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_678 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5038__B _5024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_614 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_625 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_892 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_659 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4877__B _4887_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3731__A1 _3666_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_350 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_575 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5563__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_415 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5054__A _5054_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_831 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_908 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_64 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4893__A _4893_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_676 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_613 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_624 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3302__A _3108_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_337 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4117__B _4117_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3021__B _3020_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_787 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_893 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_201 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__B1 data_out1[4] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2860__B key_in[11] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_779 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_267 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5229__A _5229_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_431 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_807 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_924 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_998 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3970__A1 _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_166 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_114 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3972__A _3972_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3420_ _3465_/A _3419_/X _3320_/X _3420_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_109_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_82 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3722__A1 _5284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_873 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_3351_ _3316_/C _3365_/B _3316_/C _3365_/B _3361_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3722__B2 _3721_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_735 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_843 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_245 VGND VPWR sky130_fd_sc_hd__decap_4
X_3282_ _3211_/X _3356_/A _3353_/A _3282_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_140_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_190 VGND VPWR sky130_fd_sc_hd__decap_6
X_5021_ _5021_/A _5019_/X _5021_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_140_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_654 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_698 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4308__A _4305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3238__B1 _3230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3212__A _3213_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_635 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3789__A1 data_in1[10] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4986__B1 _4975_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4027__B _4027_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_679 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_882 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5436__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_707 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_409 VGND VPWR sky130_fd_sc_hd__fill_2
X_4805_ _4805_/A _4815_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4738__B1 data_out2[30] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2770__B _2770_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_2997_ _2986_/A _2992_/Y _2997_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_166_239 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5139__A _5133_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4043__A _4026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_111 VGND VPWR sky130_fd_sc_hd__fill_2
X_4736_ _4699_/A _4736_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3410__B1 _3406_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_464 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3961__A1 _3908_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_306 VGND VPWR sky130_fd_sc_hd__decap_8
X_4667_ _4666_/X _4667_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4978__A _4974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_114 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3882__A _3839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_648 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_968 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_445 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5163__B1 _5052_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3618_ _3586_/A _3634_/A _3618_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_116_840 VGND VPWR sky130_fd_sc_hd__fill_2
X_4598_ _5441_/Q _4595_/B _4597_/Y _4598_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_116_862 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3713__A1 _4750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_873 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4910__B1 _5553_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_821 VGND VPWR sky130_fd_sc_hd__decap_4
X_3549_ _5154_/Y _3532_/Y _3533_/X _3534_/Y _3556_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2929__C _2989_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_692 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_757 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_898 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_375 VGND VPWR sky130_fd_sc_hd__decap_12
X_5219_ _5281_/A _5217_/X _5218_/Y _5219_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_69_470 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_941 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_45 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2945__B _2896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_676 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5321__B _5252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_827 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4218__A _4215_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_890 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_186 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_495 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4977__B1 _4997_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_860 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_713 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2961__A _2961_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_77 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_532 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4729__B1 data_out2[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_779 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_932 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_10 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_267 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5049__A _5469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_227 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3776__A1_N _2839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3401__B1 _3178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5157__A2_N _5156_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_998 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_411 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3792__A _3681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_956 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_456 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5526__RESET_B _4331_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_670 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_990 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_488 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3468__B1 _3441_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_683 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_654 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2855__B _2855_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5209__A1 _4635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4680__A2 _4674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5209__B2 _5208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_164 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4128__A _4786_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_933 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3417__B1_N _3416_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_635 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2691__B2 _2690_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3032__A _3032_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5459__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_999 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_562 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_476 VGND VPWR sky130_fd_sc_hd__fill_1
X_2920_ _2844_/Y _2920_/B _2920_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2871__A _2871_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3640__B1 _3624_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_381 VGND VPWR sky130_fd_sc_hd__decap_12
X_2851_ _2850_/A _2850_/B _2851_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_148_239 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_598 VGND VPWR sky130_fd_sc_hd__decap_4
X_5570_ _5570_/D _5129_/A _4279_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2782_ data_in2[8] _2731_/X _2733_/X _2781_/Y _5519_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_79_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4521_ _4521_/A _4577_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_615 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4798__A _5543_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_968 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5145__B1 _4572_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_659 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1019 VGND VPWR sky130_fd_sc_hd__fill_1
X_4452_ _4449_/A _4452_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_136 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_169 VGND VPWR sky130_fd_sc_hd__decap_8
X_3403_ _3400_/X _3401_/X _3402_/X _3403_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_4383_ _4397_/A _4387_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3207__A _3143_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2749__C _2749_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3171__A2 _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3334_ _3291_/A _3334_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_140_651 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_504 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_727 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_587 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_898 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_429 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_695 VGND VPWR sky130_fd_sc_hd__decap_3
X_3265_ _4639_/X _3261_/X _3262_/X _3263_/X _3264_/X _3266_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4934__A2_N _4933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1003 VGND VPWR sky130_fd_sc_hd__decap_4
X_5004_ _4985_/X _4987_/X _4978_/Y _5004_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_67_963 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2765__B _2765_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3196_ _3124_/A _3196_/B _3196_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3474__A3 _3471_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_838 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_698 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_933 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_495 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_646 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_432 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_819 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4980__B _4971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3877__A _3874_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_476 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2781__A _2852_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3575__A2_N _3574_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_830 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0_clock clkbuf_3_6_0_clock/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3596__B _3594_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_217 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_239 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_261 VGND VPWR sky130_fd_sc_hd__fill_1
X_4719_ _4718_/X _4712_/X data_out2[21] _4713_/X _4719_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_163_721 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_968 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4501__A _4501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_478 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5316__B _5281_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_915 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_68 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_79 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5151__A3 _5150_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_342 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_727 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_898 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2956__A _5222_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_183 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5332__A _5332_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4111__A1 _4096_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4111__B2 _4152_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5051__B _5038_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_944 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4147__B1_N _4146_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_977 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4890__B _4888_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_98 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_616 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3787__A _3829_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_178 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3622__B1 _3621_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_863 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_732 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5127__B1 _5116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4411__A _4411_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_927 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_618 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5226__B _5226_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_329 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_286 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3689__B1 _2689_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5142__A3 _5141_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3027__A _5527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_448 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3153__A2 _3129_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_971 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_749 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4102__A1 _3980_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3050_ _2974_/Y _3050_/B _3050_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_49_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_579 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_432 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_657 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5063__C1 _5062_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_616 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3697__A _4533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_318 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_627 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4008__D _4007_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3952_ _3915_/Y _3938_/X _3952_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_137 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2967__A2 _2965_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2903_ _4642_/A _2903_/B _2904_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_149_526 VGND VPWR sky130_fd_sc_hd__fill_2
X_3883_ _3871_/X _3878_/Y _3883_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_2834_ _2762_/Y _2795_/X _2834_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4024__C _4024_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5448__RESET_B _4424_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_209 VGND VPWR sky130_fd_sc_hd__decap_4
X_5553_ _5553_/D _5553_/Q _4299_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2765_ _5345_/B _2765_/B _2712_/X _2766_/A VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__3606__A1_N _3619_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_412 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_294 VGND VPWR sky130_fd_sc_hd__decap_3
X_4504_ _4269_/A _4504_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_172_540 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3863__C _3821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4321__A _4324_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5484_ _3677_/X _5181_/B _4381_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2696_ _2696_/A _2694_/X _2695_/Y _2696_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_133_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_478 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5136__B _5137_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_949 VGND VPWR sky130_fd_sc_hd__decap_12
X_4435_ _4438_/A _4435_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4040__B _4038_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_4366_ _4367_/A _4366_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_885 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4892__A2 _4847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_513 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2776__A _2776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_524 VGND VPWR sky130_fd_sc_hd__fill_2
X_3317_ _2885_/A _3317_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_695 VGND VPWR sky130_fd_sc_hd__decap_4
X_4297_ _4304_/A _4303_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_101_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_492 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_194 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_345 VGND VPWR sky130_fd_sc_hd__decap_12
X_3248_ _3201_/X _3248_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_132_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_451 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_900 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3447__A3 _3444_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_473 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_933 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4991__A _4992_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_389 VGND VPWR sky130_fd_sc_hd__decap_8
X_3179_ _3032_/A _3178_/A _3902_/C _3178_/Y _3180_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_82_752 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3103__C _5529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_977 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_988 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_35 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_476 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_104 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_487 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_947 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3604__B1 _3603_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_830 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_301 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3080__A1 _4638_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3080__B2 _3079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_356 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_367 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_902 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_935 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_78 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_56 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5327__A _5327_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_968 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4231__A _4231_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_938 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5046__B _5045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_757 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_245 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4885__B _4884_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_971 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_502 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_109 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4883__A2 _4872_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_684 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2686__A _4859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_299 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5062__A _4918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_602 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_911 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_270 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_793 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_465 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_999 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4406__A _4411_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2852__C _2851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5348__B1 _5324_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_879 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5541__RESET_B _4313_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_399 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4141__A _4129_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_724 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_583 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_746 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3980__A _5535_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3592__A1_N _5213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_4220_ data_in1[29] _4125_/X _4205_/X _4219_/Y _5508_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_114_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_289 VGND VPWR sky130_fd_sc_hd__decap_4
X_4151_ _3417_/X _4150_/X _3417_/X _4150_/X _4151_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_332 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_866 VGND VPWR sky130_fd_sc_hd__decap_3
X_3102_ _5355_/A _3143_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_4082_ _3299_/X _4081_/X _3299_/X _4081_/X _4082_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_505 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_676 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_782 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_229 VGND VPWR sky130_fd_sc_hd__decap_12
X_3033_ _3090_/A _3033_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_83_538 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_443 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_752 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_605 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_925 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_627 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_582 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_947 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4316__A _4312_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_295 VGND VPWR sky130_fd_sc_hd__decap_8
X_4984_ _5463_/Q _4847_/X _4942_/X _4983_/Y _5463_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3220__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_468 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3598__C1 _3597_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3935_ _5528_/Q _3935_/B _3935_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__5339__B1 _5303_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3866_ _2980_/B _3865_/X _2980_/B _3865_/X _3866_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3874__B _3852_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2817_ _5494_/Q _3012_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4011__B1 _3200_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_337 VGND VPWR sky130_fd_sc_hd__decap_4
X_3797_ _3682_/Y _3796_/X _3797_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_899 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4051__A _4050_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5536_ _3390_/X _5536_/Q _4320_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2748_ _5332_/A _2745_/X _5296_/A _2748_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_127_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_509 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_724 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_595 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_212 VGND VPWR sky130_fd_sc_hd__fill_2
X_5467_ _5035_/X _5023_/A _4401_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_746 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3890__A _3888_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_437 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3117__A2 _3115_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4418_ _4418_/A _4418_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_132_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_256 VGND VPWR sky130_fd_sc_hd__decap_12
X_5398_ _4793_/X data_out1[28] _4484_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_660 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4865__A2 _4862_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4349_ _4349_/A _4349_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_365 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_538 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_730 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3825__B1 _3815_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_752 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_56 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2953__B _2988_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_711 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_126 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_621 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3053__A1 _2973_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4135__A2_N _4134_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_66 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_321 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2800__A1 _2799_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_304 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_164 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_710 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5057__A _5028_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_540 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_724 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4896__A _4895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_470 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3305__A _3305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_505 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_376 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3024__B _3022_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4608__A2 _4605_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3816__B1 _2733_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_966 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_977 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3959__B _3936_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_465 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_947 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_593 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3040__A _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_969 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_457 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_632 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4241__B1 _4225_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_129 VGND VPWR sky130_fd_sc_hd__decap_4
X_3720_ _3701_/X _3709_/X _3681_/A _3720_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_158_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4792__A1 _4791_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4792__B2 _4782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_507 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3694__B _3692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_326 VGND VPWR sky130_fd_sc_hd__decap_8
X_3651_ _3651_/A _3649_/X _3651_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_146_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_3582_ _4537_/X _3615_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_127_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_5321_ _5252_/A _5252_/B _5321_/C _5321_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_114_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_908 VGND VPWR sky130_fd_sc_hd__decap_6
X_5252_ _5252_/A _5252_/B _5514_/Q _5252_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_88_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_716 VGND VPWR sky130_fd_sc_hd__fill_2
X_4203_ _4092_/X _4203_/B _4203_/C _4203_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_5183_ _5203_/A key_in[32] _5183_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_71 VGND VPWR sky130_fd_sc_hd__decap_12
X_4134_ _4101_/Y _4106_/X _4134_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_674 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_4065_ _4013_/Y _4064_/X _4037_/X _4065_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_37_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_763 VGND VPWR sky130_fd_sc_hd__fill_2
X_3016_ _3036_/B _3015_/X _3036_/B _3015_/X _3016_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_508 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_402 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4228__A1_N _4222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4046__A _3939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_210 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_221 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_457 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5463__RESET_B _4407_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_917 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_4967_ _4555_/A _4966_/X _4555_/A _4966_/X _4968_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3885__A _3794_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_298 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4783__A1 _4043_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3918_ _3032_/A _3917_/X _3918_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_20_630 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4783__B2 _4782_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4898_ _4908_/C _4883_/X _4873_/A _4899_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_137_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_635 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_326 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_674 VGND VPWR sky130_fd_sc_hd__fill_2
X_3849_ _3848_/X _3824_/Y _3815_/Y _3849_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_22_58 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_36 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3338__A2 key_in[120] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_829 VGND VPWR sky130_fd_sc_hd__decap_12
X_5519_ _5519_/D _2733_/C _4339_/X _5413_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_576 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_896 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_598 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5324__B _5323_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_473 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2964__A _2896_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_730 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5263__A2 _5261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3274__B2 _3273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_457 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5492__CLK _5430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_243 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_928 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_980 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4223__B1 _3395_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_963 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4774__A1 _5497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_805 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4774__B2 _4770_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2785__B1 _2761_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_838 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_624 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_623 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_337 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_696 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_668 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_122 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_540 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3019__B _3020_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_584 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_830 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_381 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_851 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4012__A2_N _4011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_351 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2858__B _2838_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_895 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5234__B key_in[34] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3035__A _3015_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_814 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_741 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5250__A _5281_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_806 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_774 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3265__A1 _4639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_519 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3265__B2 _3264_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_593 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5400__D _4796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_541 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5006__A2 _5004_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4821_ _4821_/A _4821_/B _4821_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_563 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_585 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3017__B2 _3016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_438 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_298 VGND VPWR sky130_fd_sc_hd__fill_1
X_4752_ _5229_/A _4745_/X data_out1[7] _4746_/X _4752_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3703_ _5253_/Y _5523_/Q _5514_/Q _2918_/A _3703_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_119_326 VGND VPWR sky130_fd_sc_hd__decap_12
X_4683_ _5515_/Q _4674_/X data_out2[4] _4677_/X _5406_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_88_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_605 VGND VPWR sky130_fd_sc_hd__fill_2
X_3634_ _3634_/A _3624_/X _3634_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5190__A1 _4798_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3565_ _3564_/A _3564_/B _5281_/A _3565_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_161_137 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_863 VGND VPWR sky130_fd_sc_hd__decap_3
X_5304_ _5300_/A key_in[100] _2828_/A _5304_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3740__A2 _3738_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_705 VGND VPWR sky130_fd_sc_hd__decap_12
X_3496_ _4788_/X _4794_/X _3495_/X _3496_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_102_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_598 VGND VPWR sky130_fd_sc_hd__decap_4
X_5235_ _5236_/A key_in[2] _5235_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5166_ _5165_/A _5164_/Y _5165_/X _5167_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3866__A2_N _3865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4983__B _4983_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_173 VGND VPWR sky130_fd_sc_hd__decap_12
X_4117_ _4063_/X _4117_/B _4119_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2784__A _2784_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_5097_ _5098_/A _5098_/B _5097_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5160__A _4918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_132 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3599__B _3570_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_165 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_688 VGND VPWR sky130_fd_sc_hd__decap_12
X_4048_ _3133_/A _5538_/Q _5529_/Q _4047_/Y _4048_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_140_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_582 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_766 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_703 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_216 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3008__A1 _2974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_894 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_238 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3559__A2 _3523_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4504__A _4269_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_46 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5319__B _5319_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_871 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_104 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_882 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2959__A _2959_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5335__A _5334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3192__B1 _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3731__A2 _3661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_874 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_89 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_682 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5054__B _5054_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_10 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_449 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_579 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_270 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2694__A _2695_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5070__A _5068_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_143 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5385__RESET_B _4499_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_519 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_560 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_305 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3302__B _3303_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1000 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_861 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_254 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_799 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_213 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__A1 _5287_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4414__A _4418_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__B2 _4746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_8 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_910 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__B1 _2756_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_635 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_134 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3970__A2 _3943_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5388__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3972__B _3971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_830 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2869__A _2870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5245__A _3603_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3722__A2 _5524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3350_ _3321_/Y _3349_/A _3320_/X _3419_/A _3365_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_135_1004 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_896 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_224 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_747 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_235 VGND VPWR sky130_fd_sc_hd__fill_2
X_3281_ _3217_/A _3280_/X _3241_/X _3353_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_140_877 VGND VPWR sky130_fd_sc_hd__decap_8
X_5020_ _5021_/A _5019_/X _5020_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_471 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4683__B1 data_out2[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_452 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_474 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3238__B2 _3237_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3212__B _3211_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_647 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3789__A2 _3697_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4986__A1 _4997_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_596 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_4804_ _4893_/A _4803_/Y _4805_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4738__A1 _5541_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4324__A _4324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_911 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4738__B2 _4737_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2996_ _3026_/A _2884_/B _3020_/A _2996_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__2770__C _2768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5139__B _5140_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4735_ _3493_/C _4725_/X data_out2[29] _4726_/X _5431_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4043__B _3950_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3410__A1 _4639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3410__B2 _3409_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_903 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_819 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_476 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3961__A2 _3935_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4666_ _4524_/A _4629_/D _4518_/X _4666_/D _4666_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_119_38 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4978__B _4978_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3882__B _3812_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_126 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5163__A1 _4573_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3617_ _3600_/X _3616_/Y _3634_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2779__A _2778_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4597_ _4600_/B _4597_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_162_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_619 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3713__A2 _3690_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_3548_ _5542_/Q _3548_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_351 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4910__B2 _4909_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_181 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_3479_ _3478_/X _3479_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_103_546 VGND VPWR sky130_fd_sc_hd__decap_3
X_5218_ _5192_/X _5216_/X _5218_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_57_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_920 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_5149_ _5147_/Y _5149_/B _5149_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_953 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_590 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_655 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5321__C _5321_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_839 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4218__B _4218_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_198 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_390 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4977__B2 _4976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_725 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2961__B _2961_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_900 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4234__A _4229_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4729__A1 _4728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4729__B2 _4726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_555 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3401__A1 _3325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5530__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3401__B2 _3369_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_902 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3758__A2_N _3757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_785 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_924 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_423 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_968 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5065__A _5065_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3165__B1 _3162_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_456 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4901__A1 _4900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_42 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_885 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_682 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5566__RESET_B _4284_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_419 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3468__A1 _3108_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_600 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_739 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_695 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4409__A _4411_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_441 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_452 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5209__A2 _5203_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3313__A _3170_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_603 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4128__B _4111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_422 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3032__B _3032_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_647 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_91 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2979__B1 _2974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_872 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_883 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2871__B _2871_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3640__A1 _5253_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3640__B2 _3621_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_708 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_393 VGND VPWR sky130_fd_sc_hd__decap_4
X_2850_ _2850_/A _2850_/B _2855_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4144__A _4126_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3928__C1 _3927_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_421 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _2852_/A _2779_/Y _2780_/X _2781_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_145_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_791 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3983__A _3858_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4520_ _4519_/X _4614_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_157_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_290 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4798__B _4798_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_498 VGND VPWR sky130_fd_sc_hd__decap_3
X_4451_ _4449_/A _4451_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_126 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5145__B2 _5144_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3156__B1 _3895_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3402_ _3400_/X _3401_/X _3402_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_4382_ _4381_/A _4382_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_500 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3207__B _3166_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_693 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2749__D _2748_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_833 VGND VPWR sky130_fd_sc_hd__fill_1
X_3333_ _3331_/A _3330_/X _3332_/Y _3333_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_152_490 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_663 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4105__C1 _4104_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_365 VGND VPWR sky130_fd_sc_hd__fill_2
X_3264_ _3291_/A key_in[118] _3222_/X _3264_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_39_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_611 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5202__A2_N _5201_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_29 VGND VPWR sky130_fd_sc_hd__decap_12
X_5003_ _5000_/A _4999_/X _5002_/Y _5008_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_112_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_249 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4319__A _4340_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3195_ _5013_/A _3195_/B _3195_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2765__C _2712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_806 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_975 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5403__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_658 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_444 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4959__A1 _4954_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_809 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3877__B _3876_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2781__B _2779_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5553__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_842 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4054__A _4003_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2795__B1_N _2794_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2979_ _2974_/Y _2978_/X _2974_/Y _2978_/X _2980_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_752 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3893__A _3886_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4718_ _3905_/A _4718_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_163_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_755 VGND VPWR sky130_fd_sc_hd__fill_2
X_4649_ _4577_/A _4523_/A _4649_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_123_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_408 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_46 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5332__B _5332_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4111__A2 _4109_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3133__A _3133_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_603 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_474 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_794 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_658 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_872 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_308 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3787__B _3785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3622__A1 _5514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_680 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_533 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_875 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_537 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4899__A _5552_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_251 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5127__A1 _4857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5127__B2 _4930_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_265 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4886__B1 _4885_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3689__B2 _3688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5426__CLK _5424_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_825 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_216 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4102__A2 _4098_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_430 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_709 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3043__A _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_463 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3310__B1 _3309_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3861__A1 _3750_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_625 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_422 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3978__A _4026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5576__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_978 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_230 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5063__B1 _4942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_477 VGND VPWR sky130_fd_sc_hd__decap_8
X_3951_ _3569_/A _3974_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_105 VGND VPWR sky130_fd_sc_hd__decap_6
X_2902_ _4637_/A _2898_/X _2899_/X _2900_/X _2901_/X _2903_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_31_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_853 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_3882_ _3839_/A _3812_/B _3895_/A _3882_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_52_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_2833_ _4907_/A _2830_/X _2858_/A _2838_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3377__B1 _3222_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5552_ _4549_/X _5552_/Q _4300_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4602__A _4602_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2764_ _2687_/X _2765_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_129_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_4503_ _4501_/A _4503_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_424 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4822__B1_N _4821_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_755 VGND VPWR sky130_fd_sc_hd__fill_2
X_5483_ _3653_/X _5287_/A _4382_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2695_ _2695_/A _2695_/B _2695_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_172_552 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3218__A _3145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_4434_ _4438_/A _4434_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5488__RESET_B _4377_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3130__A1_N _3125_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_118 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5417__RESET_B _4461_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4365_ _4367_/A _4365_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3316_ _3216_/A _3364_/B _3316_/C _3316_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__2776__B _2726_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_4296_ _4296_/A _4296_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4049__A _3932_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3247_ _3216_/A _3143_/B _4720_/X _3247_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_100_357 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3301__B1 _4775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_783 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_102 VGND VPWR sky130_fd_sc_hd__decap_3
X_3178_ _3178_/A _3178_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_67_794 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4991__B _4990_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5156__A2_N _5155_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_945 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3852__A1 _3875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3888__A _3770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_9 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_14 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3478__B1_N _3477_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_617 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_274 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3604__A1 _5513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_116 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_959 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_825 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_341 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_650 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3080__A2 _3076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_661 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_13 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4512__A _4515_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_593 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5327__B _5327_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4231__B _4213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3128__A _3128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_788 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_928 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5449__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5343__A _5342_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_460 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_374 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2686__B _2686_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_396 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5062__B _5060_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_506 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5293__B1 _5274_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_614 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_891 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3798__A _3682_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_786 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_650 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_323 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5348__B2 _5347_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_368 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4422__A _4422_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_700 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_891 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_744 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4141__B _4159_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_703 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3038__A _3038_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_939 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_736 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_758 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5510__RESET_B _4350_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_235 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2877__A _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5253__A _5514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3531__B1 _3408_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_514 VGND VPWR sky130_fd_sc_hd__decap_4
X_4150_ _4147_/X _4149_/B _4173_/B _4150_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_122_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_834 VGND VPWR sky130_fd_sc_hd__decap_12
X_3101_ data_in2[17] _2956_/X _3073_/X _3100_/Y _3101_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_95_344 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_569 VGND VPWR sky130_fd_sc_hd__decap_8
X_4081_ _4079_/X _4080_/X _4079_/X _4080_/X _4081_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5403__D _5403_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_666 VGND VPWR sky130_fd_sc_hd__decap_8
X_3032_ _3032_/A _3032_/B _3090_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_49_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_293 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_775 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3501__A _3501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_617 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_403 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_639 VGND VPWR sky130_fd_sc_hd__fill_2
X_4983_ _4891_/A _4983_/B _4983_/C _4983_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3220__B key_in[85] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3598__B1 _3583_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3934_ _3933_/X _3935_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_149_335 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5339__A1 _5299_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3865_ _3861_/X _3864_/Y _3865_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_31_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_379 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4332__A _4330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3874__C _3832_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2816_ _3778_/A _2819_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_3796_ _2723_/A _5527_/Q _5518_/Q _3062_/A _3796_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4011__B2 _4010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_530 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_744 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_27 VGND VPWR sky130_fd_sc_hd__decap_3
X_2747_ _5325_/A _5332_/A _2746_/Y _2749_/C VGND VPWR sky130_fd_sc_hd__o21a_4
X_5535_ _3363_/X _5535_/Q _4321_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_511 VGND VPWR sky130_fd_sc_hd__decap_8
X_5466_ _5022_/Y _5013_/A _4402_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3890__B _3889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_544 VGND VPWR sky130_fd_sc_hd__decap_8
X_4417_ _4418_/A _4417_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_555 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2787__A _2898_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5397_ _4792_/X data_out1[27] _4485_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_132_268 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3522__B1 _3510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_983 VGND VPWR sky130_fd_sc_hd__fill_1
X_4348_ _4349_/A _4348_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_834 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3084__A1_N _3128_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_845 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_867 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_4279_ _4276_/X _4279_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_28_901 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_699 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3286__C1 _3285_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_282 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3825__B2 _3824_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_742 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2721__A2_N _2720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_455 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4507__A _4504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_572 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3053__A2 _3006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_633 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_300 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_56 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_834 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_132 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_78 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2800__A2 _2799_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5338__A _2707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_867 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_816 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_891 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_337 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5057__B _5057_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3355__B1_N _3354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_850 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_736 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_554 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3305__B _3305_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_86 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_804 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_997 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3024__C _3023_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_325 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3816__A1 _2735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3816__B2 _3075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_30 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_347 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3605__A1_N _5242_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4417__A _4418_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_764 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3959__C _3912_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_252 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3321__A _3320_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_712 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_296 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_745 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3040__B key_in[48] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_611 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4241__A1 _3395_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_644 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4792__A2 _4781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_299 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5248__A _5246_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_828 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4152__A _4152_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3650_ _3651_/A _3649_/X _3650_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_9_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_349 VGND VPWR sky130_fd_sc_hd__decap_8
X_3581_ _5222_/A _3581_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_155_872 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3991__A _4775_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5320_ data_in2[4] _5222_/X _5283_/X _5319_/X _5515_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_127_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_725 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_393 VGND VPWR sky130_fd_sc_hd__decap_4
X_5251_ data_in2[2] _5222_/X _5224_/X _5250_/X _5513_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_114_235 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_4202_ _4195_/X _4232_/C _4203_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3504__B1 _3502_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_780 VGND VPWR sky130_fd_sc_hd__decap_12
X_5182_ _3578_/A _3671_/A _5181_/X _5182_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_96_642 VGND VPWR sky130_fd_sc_hd__decap_4
X_4133_ _4000_/Y _4131_/X _4132_/X _4133_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_110_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_141 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_837 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_997 VGND VPWR sky130_fd_sc_hd__fill_2
X_4064_ _4778_/X _4036_/X _4064_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_56_539 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_3015_ _3015_/A _2966_/X _3015_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_83_358 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4327__A _4330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3231__A _3231_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_786 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_263 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4046__B _4045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_929 VGND VPWR sky130_fd_sc_hd__decap_12
X_4966_ _4921_/X _4965_/X _4966_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_110 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3885__B _3884_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_132 VGND VPWR sky130_fd_sc_hd__decap_4
X_3917_ _3904_/X _3915_/Y _3916_/X _3917_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__4783__A2 _4781_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4897_ _5456_/Q _4900_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5158__A _5159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_3848_ _3587_/B _3848_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5432__RESET_B _4443_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4997__A _4555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_541 VGND VPWR sky130_fd_sc_hd__fill_2
X_3779_ _3778_/X _3780_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_861 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_319 VGND VPWR sky130_fd_sc_hd__fill_2
X_5518_ _5518_/D _5518_/Q _4341_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_382 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_224 VGND VPWR sky130_fd_sc_hd__decap_12
X_5449_ _4826_/X _4817_/A _4423_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_706 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_36 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3406__A _3337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_333 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_249 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_804 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_986 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_325 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2964__B _2964_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_904 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_915 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3141__A _3170_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_274 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_33 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_44 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2980__A _2980_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3591__A1_N _3573_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_469 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_789 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4038__B1_N _4037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4223__B2 _3521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_439 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_17 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_299 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_975 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4774__A2 _4769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_986 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2785__A1 _2762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5068__A _5068_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_102 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_635 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4700__A _4700_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_691 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_842 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_clock clkbuf_3_6_0_clock/A clkbuf_3_7_0_clock/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_152_853 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_363 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3316__A _3216_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_717 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_897 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_620 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3035__B _3014_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_249 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_750 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5239__B1 _4817_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5250__B _5278_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_347 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_689 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3265__A2 _3261_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3051__A _2977_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4820_ _4541_/A _4819_/X _4541_/A _4819_/X _4821_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_929 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4214__A1 _4794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_428 VGND VPWR sky130_fd_sc_hd__decap_4
X_4751_ _4750_/X _4745_/X data_out1[6] _4746_/X _4751_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_105_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_474 VGND VPWR sky130_fd_sc_hd__fill_2
X_3702_ _3681_/A _3701_/X _3702_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_4682_ _5514_/Q _4674_/X data_out2[3] _4677_/X _4682_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_119_338 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_658 VGND VPWR sky130_fd_sc_hd__decap_12
X_3633_ _3615_/A _3570_/B _5287_/A _3633_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_146_168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_872 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4610__A _4609_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3564_ _3564_/A _3564_/B _3564_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__5190__A2 _5189_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5303_ _5303_/A _2828_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_3495_ _3178_/Y _3495_/B _3495_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_103_717 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_897 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3226__A _5468_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_694 VGND VPWR sky130_fd_sc_hd__decap_8
X_5234_ _5234_/A key_in[34] _5234_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_102_227 VGND VPWR sky130_fd_sc_hd__fill_1
X_5165_ _5165_/A _5164_/Y _5165_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_506 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4983__C _4983_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1005 VGND VPWR sky130_fd_sc_hd__fill_2
X_4116_ _4784_/X _4083_/X _4115_/X _4120_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_83_100 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_483 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_794 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2784__B _2779_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5096_ _5081_/X _5096_/B _5098_/B VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_56_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_185 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5160__B _5160_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3599__C _5481_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4047_ _5538_/Q _4047_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_37_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_701 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_594 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3896__A _3895_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_907 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_778 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_406 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3008__A2 _2978_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_228 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1000 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_239 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_299 VGND VPWR sky130_fd_sc_hd__decap_12
X_4949_ _4949_/A _4949_/B _4949_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_165_400 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3964__B1 _3131_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5319__C _5319_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_483 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_116 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4520__A _4519_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_691 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5335__B _5309_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3192__A1 _3145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_672 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3136__A _3073_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_800 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_951 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2975__A _2913_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_984 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5351__A _5351_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_794 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2694__B _2695_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_645 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_61 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5070__B _5067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_509 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5501__D _4070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_372 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_299 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__A2 _4745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_64 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_772 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_247 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__A1 _4637_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_794 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_86 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__B2 _2757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_922 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_647 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_669 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_454 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_639 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4430__A _4426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_127 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2869__B _2870_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5245__B _5245_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_715 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4227__A1_N _3535_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_3280_ _4718_/X _3280_/B _3280_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_124_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_940 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2885__A _2885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4683__A1 _5515_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5261__A _5261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_910 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4683__B2 _4677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_678 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5411__D _5411_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_497 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3498__A1_N _3496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_594 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_659 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4986__A2 _4976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_851 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4605__A _4646_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_748 VGND VPWR sky130_fd_sc_hd__decap_12
X_4803_ _4656_/X _4803_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4738__A2 _4736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3421__A1_N _3436_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2995_ data_in2[14] _2956_/X _2958_/X _2994_/Y _5525_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__2770__D _2769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_400 VGND VPWR sky130_fd_sc_hd__decap_12
X_4734_ _5540_/Q _3493_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_159_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_293 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4043__C _4043_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3410__A2 _3404_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4665_ _4664_/X _3676_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_135_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_639 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3882__C _3895_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4340__A _4340_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3616_ _3606_/X _3616_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5163__A2 _5155_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4596_ _4595_/X _4600_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_661 VGND VPWR sky130_fd_sc_hd__decap_8
X_3547_ _3521_/X _3537_/X _3545_/B _3564_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_116_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2692__A1_N _5356_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_300 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_171 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5482__CLK _5456_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_49 VGND VPWR sky130_fd_sc_hd__fill_2
X_3478_ _3475_/X _3477_/B _3477_/X _3478_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_88_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_193 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5320__C1 _5319_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5217_ _5192_/X _5216_/X _5217_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_15 VGND VPWR sky130_fd_sc_hd__decap_3
X_5148_ _5132_/Y _5148_/B _5149_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2685__B1 _5368_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_580 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_5079_ _4566_/A _5078_/X _4566_/A _5078_/X _5079_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4515__A _4515_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_586 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4011__A2_N _4010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_748 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4729__A2 _4725_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4234__B _4234_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_63 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_731 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3401__A2 _3370_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_989 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_414 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4250__A _4577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_959 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_842 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5065__B _5051_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3165__B2 _3164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_864 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4901__A2 _4899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_897 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_269 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_910 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3468__A2 _3251_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5081__A _5080_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_932 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_291 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3313__B _3313_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_818 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5209__A3 _5204_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_924 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_434 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5535__RESET_B _4321_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3850__A2_N _3849_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_309 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2979__B2 _2978_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4425__A _4422_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_350 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_501 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3640__A2 _2735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4144__B _4090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4151__A1_N _3417_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_720 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3928__B1 _3902_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2780_ _2778_/A _2777_/X _2780_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_589 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_753 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3983__B _3981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_786 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5256__A _5256_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_105 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4160__A _4788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_796 VGND VPWR sky130_fd_sc_hd__decap_8
X_4450_ _4449_/A _4450_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_172_745 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3156__A1 _3012_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3401_ _3325_/X _3370_/X _3332_/Y _3178_/Y _3369_/X _3401_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__3156__B2 _3155_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4381_ _4381_/A _4381_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5406__D _5406_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_661 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_992 VGND VPWR sky130_fd_sc_hd__fill_2
X_3332_ _3331_/X _3332_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_140_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_867 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4105__B1 _4078_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_567 VGND VPWR sky130_fd_sc_hd__fill_1
X_3263_ _3293_/A key_in[86] _3263_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_58_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_675 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_910 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3803__A2_N _3802_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5002_ _5001_/X _5002_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3194_ _5023_/A _3228_/B _5023_/A _3228_/B _3199_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_280 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_604 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_166 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4959__A2 _4958_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_979 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_456 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4335__A _4339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3092__B1 _3937_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2781__C _2780_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_821 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3990__A1_N _3987_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_854 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4054__B _4031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_38 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3919__B1 _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_589 VGND VPWR sky130_fd_sc_hd__decap_12
X_2978_ _2912_/X _2975_/X _2977_/Y _2978_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3893__B _3892_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_241 VGND VPWR sky130_fd_sc_hd__decap_3
X_4717_ _3175_/A _4712_/X data_out2[20] _4713_/X _5422_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4592__B1 _4591_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_745 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_436 VGND VPWR sky130_fd_sc_hd__fill_2
X_4648_ _4645_/X _4671_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_907 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_458 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_929 VGND VPWR sky130_fd_sc_hd__fill_2
X_4579_ _4579_/A _5256_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_150_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_534 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_664 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4647__A1 _4256_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_910 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_36 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3414__A _3342_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_58 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3133__B _3133_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_453 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_762 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_615 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_486 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_6_0_clock clkbuf_4_7_0_clock/A _5424_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_73_957 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_283 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_840 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5378__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_361 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3083__B1 _3048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3622__A2 _2733_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_821 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_383 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_832 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_692 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_22 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2830__B1 _2826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_539 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_731 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4899__B _4899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_99 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3386__A1 _4728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5076__A _5076_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5127__A2 _5125_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_907 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_277 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4886__A1 _4885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_276 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_504 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3324__A _3155_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_537 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_932 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_943 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_442 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_751 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3310__A1 _3287_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3861__A2 _3859_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3978__B _3950_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5063__A1 _5469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_242 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_873 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4155__A _3396_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3950_ _3839_/A _3950_/B _5497_/Q _3950_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_63_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_361 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_832 VGND VPWR sky130_fd_sc_hd__fill_2
X_2901_ _2898_/A key_in[108] _2828_/A _2901_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__2821__B1 _2799_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3881_ data_in1[14] _3837_/X _3857_/X _3880_/Y _5493_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3994__A _3979_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_865 VGND VPWR sky130_fd_sc_hd__decap_12
X_2832_ _2832_/A _2858_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3377__A1 _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_904 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_550 VGND VPWR sky130_fd_sc_hd__fill_2
X_5551_ _4548_/X _4908_/C _4301_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2763_ _2686_/Y _2711_/Y _2770_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_145_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_274 VGND VPWR sky130_fd_sc_hd__decap_12
X_4502_ _4501_/A _4502_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_745 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_2694_ _2695_/A _2695_/B _2694_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_5482_ _3632_/X _5260_/A _4384_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_144_233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_778 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3218__B key_in[53] VGND VPWR sky130_fd_sc_hd__diode_2
X_4433_ _4419_/A _4438_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_810 VGND VPWR sky130_fd_sc_hd__decap_12
X_4364_ _4367_/A _4364_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3315_ _5355_/A _3364_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_375 VGND VPWR sky130_fd_sc_hd__decap_12
X_4295_ _4296_/A _4295_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3234__A _3233_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_314 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_483 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5457__RESET_B _4414_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3246_ data_in2[21] _3172_/X _3216_/X _3245_/Y _5532_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4049__B _4048_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3301__A1 _3158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_369 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5520__CLK _5402_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3301__B2 _3466_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3177_ _4582_/X _3176_/X _3177_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_39_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3852__A2 _3850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_423 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3888__B _3887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_136 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_15 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_927 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_37 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_938 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_48 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3604__A2 _5518_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4058__A1_N _4046_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_837 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3080__A3 _3077_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_325 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_504 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_386 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_548 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_211 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_436 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3128__B _3128_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_406 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_981 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_515 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3144__A _3144_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_19 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5062__C _5061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5293__A1 _3626_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5293__B2 _5262_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4959__B1_N _4958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_710 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_626 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3798__B _3796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_968 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_456 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_681 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2803__B1 _2796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_353 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4703__A _5524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_172 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_357 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_723 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3319__A _3465_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_520 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3038__B _3037_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_970 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5216__A2_N _5215_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_225 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_439 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2877__B _2876_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_962 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3531__A1 _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5543__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_601 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3054__A _2975_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3100_ _2927_/A _3098_/Y _3099_/X _3100_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_122_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_846 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5550__RESET_B _4302_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4080_ _4052_/X _4055_/Y _4050_/X _4080_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_95_356 VGND VPWR sky130_fd_sc_hd__fill_2
X_3031_ _2714_/Y _3030_/A _2714_/A _3233_/A _3032_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_95_367 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2893__A _2872_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3295__B1 _3293_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_957 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_467 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3501__B key_in[29] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_275 VGND VPWR sky130_fd_sc_hd__fill_2
X_4982_ _4982_/A _4980_/X _4983_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_17_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_990 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_437 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3598__A1 data_in1[1] VGND VPWR sky130_fd_sc_hd__diode_2
X_3933_ _3721_/Y _4720_/X _2989_/A _3932_/Y _3933_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4795__B1 data_out1[29] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_651 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_971 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5339__A2 key_in[101] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_347 VGND VPWR sky130_fd_sc_hd__decap_12
X_3864_ _3843_/Y _3862_/Y _3863_/Y _3864_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_20_835 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_306 VGND VPWR sky130_fd_sc_hd__decap_4
X_2815_ _5358_/A _2814_/X _2815_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_164_317 VGND VPWR sky130_fd_sc_hd__decap_8
X_3795_ _3773_/X _3774_/X _3819_/A _3795_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3229__A _3228_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_891 VGND VPWR sky130_fd_sc_hd__decap_12
X_5534_ _3314_/X _5534_/Q _4322_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_157_391 VGND VPWR sky130_fd_sc_hd__fill_2
X_2746_ _2745_/X _2746_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_145_542 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_704 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_715 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_789 VGND VPWR sky130_fd_sc_hd__fill_2
X_5465_ _5012_/X _4996_/A _4403_/X _5579_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_4416_ _4418_/A _4416_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5396_ _4790_/X data_out1[26] _4486_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2787__B key_in[41] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3522__A1 _4661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_504 VGND VPWR sky130_fd_sc_hd__fill_2
X_4347_ _4340_/A _4349_/A VGND VPWR sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0_clock clkbuf_0_clock/X clkbuf_2_3_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__2730__C1 _2729_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_345 VGND VPWR sky130_fd_sc_hd__decap_12
X_4278_ _4276_/X _4278_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_101_656 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3899__A _3883_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_507 VGND VPWR sky130_fd_sc_hd__decap_4
X_3229_ _3228_/X _3199_/Y _3229_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_86_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_710 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3286__B1 _3247_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_776 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_618 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_798 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_768 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_640 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1004 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_779 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_662 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_13 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_982 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4523__A _4523_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_684 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5416__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_667 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_846 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5338__B key_in[69] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_306 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3139__A _3139_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_862 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_553 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_350 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5566__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_895 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_748 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5379__RESET_B _4506_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_544 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_578 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_150 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5504__D _4143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_902 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_827 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3816__A2 _5528_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_743 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5018__A1 _5017_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_clock clkbuf_3_2_0_clock/A clkbuf_4_7_0_clock/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_93_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_437 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4777__B1 data_out1[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_623 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4241__A2 _3521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_971 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4433__A _4419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_161 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_807 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_132 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5248__B _5249_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_166 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4152__B _4136_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_198 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3201__B1 _3188_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3580_ data_in1[0] _3391_/X _3570_/X _3579_/X _3580_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_155_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_850 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3991__B _3990_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_704 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2888__A _2999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_512 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_371 VGND VPWR sky130_fd_sc_hd__fill_1
X_5250_ _5281_/A _5278_/B _5250_/C _5250_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_47_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_258 VGND VPWR sky130_fd_sc_hd__fill_2
X_4201_ _4195_/X _4232_/C _4203_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3504__A1 _4640_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_813 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3504__B2 _3503_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5414__D _5414_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_824 VGND VPWR sky130_fd_sc_hd__fill_2
X_5181_ _3577_/A _5181_/B _5181_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_123_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_40 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_846 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_62 VGND VPWR sky130_fd_sc_hd__fill_2
X_4132_ _4000_/Y _4131_/X _4132_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3400__B1_N _3399_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_95 VGND VPWR sky130_fd_sc_hd__decap_6
X_4063_ _4014_/X _4038_/X _4063_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_3_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3268__B1 _3267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_710 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_592 VGND VPWR sky130_fd_sc_hd__fill_2
X_3014_ _3014_/A _3014_/B _3036_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_25_905 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_798 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_735 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5439__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4768__B1 data_out1[15] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_4965_ _4554_/A _4955_/X _4965_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4343__A _4341_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3916_ _3904_/X _3915_/Y _3916_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4896_ _4895_/X _4896_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_149_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_604 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2983__A1_N _2998_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5158__B _5159_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_3847_ _2939_/X _3846_/X _2939_/X _3846_/X _3847_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_648 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_147 VGND VPWR sky130_fd_sc_hd__decap_6
X_3778_ _3778_/A _3777_/X _3778_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4997__B _4965_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5517_ _5517_/D _5517_/Q _4342_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_106_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_2729_ _2852_/A _2727_/X _2728_/Y _2729_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_161_810 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_737 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5174__A _2885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_180 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_394 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5472__RESET_B _4395_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5448_ _4816_/X _5448_/Q _4424_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_887 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_718 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_589 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3406__B key_in[90] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5401__RESET_B _4480_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5379_ _4755_/X data_out1[9] _4506_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_345 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_816 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_453 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_209 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_827 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4518__A _4518_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2964__C _2895_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3422__A _3395_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_186 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_220 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3141__B _3139_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_927 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_415 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5233__A1_N _5231_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_286 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_757 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4759__B1 data_out1[10] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2980__B _2980_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_960 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__A _4524_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_954 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_621 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_790 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_998 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2785__A2 _2770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_829 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_120 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5068__B _5067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_647 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_564 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4931__B1 _2907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_117 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_128 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5084__A _5084_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_865 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_875 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3316__B _3364_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3498__B1 _3496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_363 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_654 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5239__B2 _5238_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_762 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4428__A _4426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_635 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3332__A _3331_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5250__C _5250_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_540 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3265__A3 _3262_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3051__B _3050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_735 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_521 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_768 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4214__A2 _4212_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4163__A _4158_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4750_ _5200_/A _4750_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_159_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1013 VGND VPWR sky130_fd_sc_hd__decap_6
X_3701_ _3680_/X _3689_/Y _3701_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_615 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_963 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_306 VGND VPWR sky130_fd_sc_hd__decap_6
X_4681_ _5513_/Q _4674_/X data_out2[2] _4677_/X _4681_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_147_626 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5409__D _4690_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_3632_ data_in1[3] _3581_/X _3615_/X _3631_/X _3632_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_127_350 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_629 VGND VPWR sky130_fd_sc_hd__fill_1
X_3563_ _3557_/X _3562_/X _3557_/X _3562_/X _3564_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_692 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3507__A _3505_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2720__A2_N _2719_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5302_ _5301_/A key_in[68] _5302_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_154_191 VGND VPWR sky130_fd_sc_hd__decap_6
X_3494_ _3465_/B _3480_/Y _3465_/A _3510_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3226__B _3226_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_375 VGND VPWR sky130_fd_sc_hd__fill_2
X_5233_ _5231_/Y _5258_/A _5231_/Y _5258_/A _5233_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_386 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4150__A1 _4147_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5164_ _5478_/Q _5164_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_96_440 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_518 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_602 VGND VPWR sky130_fd_sc_hd__decap_12
X_4115_ _4115_/A _4115_/B _4115_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_56_304 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4338__A _4339_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5095_ _5090_/Y _5093_/X _5109_/B _5098_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_56_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5160__C _5160_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4046_ _3939_/X _4045_/X _4046_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_17_38 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_329 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_830 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3896__B _3894_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5169__A _5169_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_229 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_727 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4073__A _3939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1012 VGND VPWR sky130_fd_sc_hd__decap_8
X_4948_ _4943_/Y _4946_/X _4947_/X _4951_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_149_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3964__B2 _3963_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_412 VGND VPWR sky130_fd_sc_hd__decap_8
X_4879_ _4877_/X _4878_/X _4879_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_21_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_445 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4801__A _4656_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_456 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_489 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4913__B1 _4885_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_128 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_320 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3192__A2 key_in[116] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_138 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_353 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3136__B _3096_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_589 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_397 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_537 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_941 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2975__B _2938_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_153 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5351__B _5351_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_849 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2875__A1_N _2857_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_657 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_540 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3101__C1 _3100_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_616 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2991__A _2988_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_768 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_267 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_384 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__A2 _2754_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_784 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_934 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_283 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5157__B1 _5154_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5394__RESET_B _4488_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_467 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_607 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_180 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_876 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_662 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_364 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_727 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_194 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_952 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4683__A2 _4674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_922 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_933 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3062__A _3062_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_977 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3997__A _4026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_532 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_148 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A clkbuf_2_0_0_clock/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__4605__B _4605_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_4802_ _4857_/A _4802_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_21_204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_395 VGND VPWR sky130_fd_sc_hd__decap_12
X_2994_ _2927_/A _2992_/Y _2993_/X _2994_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_15_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_209 VGND VPWR sky130_fd_sc_hd__fill_1
X_4733_ _5539_/Q _4725_/X data_out2[28] _4726_/X _4733_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_147_412 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3410__A3 _3405_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_18 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4621__A _5301_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4664_ _3584_/B _4664_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_629 VGND VPWR sky130_fd_sc_hd__fill_1
X_3615_ _3615_/A _3570_/B _5260_/A _3615_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4595_ _5441_/Q _4595_/B _4595_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3418__A2_N _3417_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_640 VGND VPWR sky130_fd_sc_hd__fill_2
X_3546_ data_in2[30] _3391_/X _3519_/X _3545_/X _3546_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_116_865 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_526 VGND VPWR sky130_fd_sc_hd__decap_12
X_3477_ _3475_/X _3477_/B _3477_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_345 VGND VPWR sky130_fd_sc_hd__decap_8
X_5216_ _4679_/X _5215_/X _4679_/X _5215_/X _5216_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5320__B1 _5283_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_440 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_782 VGND VPWR sky130_fd_sc_hd__fill_2
X_5147_ _5143_/X _5145_/Y _5146_/X _5147_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XANTENNA__4068__A _4068_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_410 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2685__A1 _4636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2685__B2 _5369_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_966 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_49 VGND VPWR sky130_fd_sc_hd__fill_2
X_5078_ _5037_/X _5077_/X _5078_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_57_679 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2689__A2_N _2688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_178 VGND VPWR sky130_fd_sc_hd__decap_8
X_4029_ _3905_/Y _4028_/X _4029_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_25_521 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_690 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3700__A _3569_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_660 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_69 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_598 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_215 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3401__A3 _3332_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_220 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4531__A _4546_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3861__B1_N _3860_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_607 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_798 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_403 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_clock clkbuf_4_3_0_clock/A _5382_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__4250__B _4578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_681 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_139 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3147__A _3077_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_191 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_876 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2986__A _2986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5311__B1 _5310_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_664 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_922 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5512__D _5220_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3873__B1 _3872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_668 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3313__C _3312_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_914 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5075__C1 _5074_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_882 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_532 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_446 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_468 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_513 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5575__RESET_B _4272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4144__C _3231_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1002 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3928__A1 data_in1[16] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5504__RESET_B _4357_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4441__A _4443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_765 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5256__B _5256_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4160__B _4137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_448 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3057__A _3051_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3400_ _3396_/X _3398_/X _3399_/X _3400_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3156__A2 _3155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_4380_ _4381_/A _4380_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_4_970 VGND VPWR sky130_fd_sc_hd__fill_2
X_3331_ _3331_/A _3330_/X _3331_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_113_824 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2896__A _2896_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4105__A1 _4051_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3262_ _3293_/A key_in[22] _3262_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_140_687 VGND VPWR sky130_fd_sc_hd__decap_8
X_5001_ _5001_/A _5001_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5422__D _5422_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5079__A1_N _4566_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3193_ _4638_/X _3189_/X _3190_/X _3191_/X _3192_/X _3228_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_67_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_443 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_616 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_649 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4616__A _4615_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3520__A _5541_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_468 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3092__B2 _3091_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5369__B1 _2828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4054__C _4008_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_866 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3919__A1 _3032_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2977_ _2905_/A _2976_/X _2937_/X _2977_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4716_ _3143_/C _4712_/X data_out2[19] _4713_/X _5421_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4592__A1 _4589_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4351__A _4349_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_927 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_4647_ _4256_/A _4645_/X _4646_/X _5435_/D VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3987__A2_N _3986_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_907 VGND VPWR sky130_fd_sc_hd__decap_8
X_4578_ _4578_/A _5172_/A _4579_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_2_918 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_418 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_982 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_417 VGND VPWR sky130_fd_sc_hd__fill_2
X_3529_ _3529_/A key_in[30] _3529_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_1_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_632 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_194 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_568 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4647__A2 _4645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_698 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3414__B _3414_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_281 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4211__A1_N _3508_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_627 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_936 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4526__A _4650_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3607__B1 _3601_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3430__A _3431_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3083__A1 _3128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2830__A1 _4637_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2830__B2 _2829_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_899 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5357__A _5323_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_398 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3386__A2 _3385_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4261__A _4629_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_712 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_286 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5127__A3 _5126_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_437 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5507__D _4204_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_919 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_789 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4886__A2 _4884_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_610 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_71 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2897__A1 _2896_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5092__A _5052_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_985 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_516 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3324__B _3324_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3846__B1 _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_977 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3310__A2 _3309_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_785 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_733 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3978__C _4775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4436__A _4438_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3753__B1_N _3752_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3340__A _5076_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_446 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5063__A2 _4995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4155__B _4154_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_671 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_896 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_822 VGND VPWR sky130_fd_sc_hd__fill_2
X_2900_ _2790_/A key_in[76] _2900_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2691__A1_N _5358_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_3880_ _3835_/A _3878_/Y _3879_/X _3880_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__2821__A1 _2741_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5472__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2821__B2 _2799_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3994__B _4015_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_877 VGND VPWR sky130_fd_sc_hd__decap_8
X_2831_ _4907_/A _2830_/X _2832_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_387 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5267__A _5236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5220__C1 _5219_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_540 VGND VPWR sky130_fd_sc_hd__decap_4
X_5550_ _5550_/D _4874_/A _4302_/X _5547_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3377__A2 key_in[121] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4171__A _4073_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2762_ _4882_/A _2759_/B _2761_/Y _2762_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_129_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4501_ _4501_/A _4501_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_521 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_286 VGND VPWR sky130_fd_sc_hd__decap_8
X_5481_ _3614_/X _5481_/Q _4385_/X _5456_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5417__D _4708_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2693_ _5321_/C _5348_/X _5351_/X _2695_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_117_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_245 VGND VPWR sky130_fd_sc_hd__decap_4
X_4432_ _4426_/X _4432_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_822 VGND VPWR sky130_fd_sc_hd__decap_12
X_4363_ _4367_/A _4363_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_153_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_941 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3515__A _3516_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_3314_ data_in2[23] _3172_/X _3287_/X _3313_/Y _3314_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_99_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_4294_ _4296_/A _4294_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_676 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3234__B _3233_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_538 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_838 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_326 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_186 VGND VPWR sky130_fd_sc_hd__fill_2
X_3245_ _3170_/A _3245_/B _3244_/X _3245_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_100_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_741 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3301__A2 _3300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2962__B1_N _3015_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3176_ _3060_/B _3176_/B _3162_/X _3163_/X _3176_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_27_605 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_774 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4346__A _4341_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5497__RESET_B _4366_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_593 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_435 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3250__A _4582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_232 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5426__RESET_B _4451_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_788 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_298 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_855 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_674 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_516 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4014__B1 _4013_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5177__A _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3128__C _3057_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_610 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_930 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5212__B1_N _5211_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_131 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_996 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_527 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3144__B _3139_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_495 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5293__A2 _5292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_722 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4256__A _4256_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3160__A _3160_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5495__CLK _5429_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2803__B2 _2802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_866 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5087__A _5087_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_713 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3764__C1 _3763_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3319__B _3319_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_381 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_716 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_575 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_597 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3335__A _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3531__A2 key_in[126] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_313 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3054__B _3050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_280 VGND VPWR sky130_fd_sc_hd__decap_12
X_3030_ _3030_/A _3233_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_37_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_379 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3295__A1 _4639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2893__B _2871_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_402 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3295__B2 _3294_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_785 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_936 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_435 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_530 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3070__A _3069_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_574 VGND VPWR sky130_fd_sc_hd__fill_2
X_4981_ _4982_/A _4980_/X _4983_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_17_693 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4795__A1 _4794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_449 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3598__A2 _3581_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3932_ _4720_/A _3932_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4795__B2 _4677_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_663 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_326 VGND VPWR sky130_fd_sc_hd__fill_2
X_3863_ _3818_/X _3844_/X _3821_/Y _3863_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_20_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_359 VGND VPWR sky130_fd_sc_hd__decap_6
X_2814_ _2702_/X _2722_/B _2813_/Y _2814_/D _2814_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_31_184 VGND VPWR sky130_fd_sc_hd__decap_3
X_3794_ _3794_/A _3793_/X _3794_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3229__B _3199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_5533_ _3286_/X _4720_/A _4323_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2745_ _2744_/X _2745_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_768 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_554 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_5464_ _5464_/D _5464_/Q _4406_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_172_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_4415_ _4418_/A _4415_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5395_ _5395_/D data_out1[25] _4487_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3245__A _3170_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_4346_ _4341_/A _4346_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3522__A2 _3510_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_302 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2730__B1 _2698_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_484 VGND VPWR sky130_fd_sc_hd__decap_4
X_4277_ _4276_/X _4277_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_86_357 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3899__B _3921_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_668 VGND VPWR sky130_fd_sc_hd__decap_3
X_3228_ _5023_/A _3228_/B _3228_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3286__A1 data_in2[22] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_880 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_733 VGND VPWR sky130_fd_sc_hd__fill_2
X_3159_ _3182_/B _3159_/B _3183_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_70_703 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_788 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4804__A _4893_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1016 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_994 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_25 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_471 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_313 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_679 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_702 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_829 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_178 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4532__A2_N _4531_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3139__B _3138_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_841 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3155__A _3155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_952 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_825 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2721__B1 _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2994__A _2927_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5166__B1_N _5165_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_977 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_519 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_50 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_593 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5520__D _2811_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_446 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5018__A2 _5017_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_703 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4777__A1 _3010_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_630 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4777__B2 _4770_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2807__B1_N _2806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_983 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_668 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_880 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5510__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3201__B2 _3200_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_840 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3756__A2_N _3755_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_885 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2888__B _2887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_373 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2960__B1 _3778_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_895 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_749 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3065__A _3065_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4200_ _4178_/X _4196_/Y _4200_/C _4200_/D _4232_/C VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__3504__A2 _3500_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4057__A1_N _3273_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5180_ _5327_/A _3671_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_122_270 VGND VPWR sky130_fd_sc_hd__decap_4
X_4131_ _3905_/Y _5541_/Q _4718_/X _3520_/Y _4131_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_110_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_933 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5280__A _5277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_666 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_508 VGND VPWR sky130_fd_sc_hd__decap_8
X_4062_ _4043_/C _4058_/X _4115_/A _4068_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3268__A1 _5469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_3013_ _3012_/A _3012_/B _3014_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5430__D _4733_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_243 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_980 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_427 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_449 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4768__A1 _3895_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4768__B2 _4758_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4624__A _3077_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4964_ _5462_/Q _3052_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3709__A2_N _3708_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3915_ _3058_/X _3914_/X _3058_/X _3914_/X _3915_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_149_123 VGND VPWR sky130_fd_sc_hd__decap_3
X_4895_ _5223_/A _4918_/A _4895_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_32_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_808 VGND VPWR sky130_fd_sc_hd__decap_3
X_3846_ _3844_/X _3845_/X _3844_/X _3845_/X _3846_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_627 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_104 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_178 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_329 VGND VPWR sky130_fd_sc_hd__fill_2
X_3777_ _3768_/Y _3776_/X _3768_/Y _3776_/X _3777_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4997__C _4997_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2728_ _2728_/A _2728_/B _2728_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_5516_ _5354_/X _5516_/Q _4343_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_106_727 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_833 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_844 VGND VPWR sky130_fd_sc_hd__decap_8
X_5447_ _4807_/X _4798_/B _4425_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_106_749 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_365 VGND VPWR sky130_fd_sc_hd__decap_4
X_5378_ _4753_/X data_out1[8] _4507_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_460 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_782 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_4329_ _4330_/A _4329_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_493 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_121 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_644 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_465 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_700 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5441__RESET_B _4432_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_379 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_839 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3422__B _3421_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3141__C _3141_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_872 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4208__B1 _4207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4759__A1 _3778_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5215__A2_N _5226_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4534__A _4533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_544 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4759__B2 _4758_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_79 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_972 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_994 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__B _4629_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_432 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_611 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5533__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_977 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_666 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_103 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2989__A _2989_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_841 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_659 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_863 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_158 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4931__A1 _4870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4931__B2 _4930_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5515__D _5515_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_65 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3316__C _3316_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5529__RESET_B _4328_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_771 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4695__B1 data_out2[10] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3498__B2 _3497_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_666 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3613__A _3579_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_799 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_533 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4444__A _4443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_950 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_410 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4163__B _4163_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_994 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_780 VGND VPWR sky130_fd_sc_hd__fill_2
X_3700_ _3569_/A _3788_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4680_ _4679_/X _4674_/X data_out2[1] _4677_/X _5403_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_169_90 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3631_ _3579_/A _3631_/B _3630_/Y _3631_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__2899__A _2790_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5275__A _5256_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3562_ _3562_/A _3562_/B _3562_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_143_822 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_513 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_5301_ _5301_/A key_in[4] _5301_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_310 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3507__B _3507_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_855 VGND VPWR sky130_fd_sc_hd__decap_8
X_3493_ _3519_/A _3364_/B _3493_/C _3493_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__5425__D _5425_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_5232_ _5199_/Y _5361_/A _5181_/X _5201_/X _5258_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_5163_ _4573_/A _5155_/X _5052_/A _5167_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4150__A2 _4149_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_953 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2697__C1 _2696_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4619__A _5236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3523__A _3368_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_975 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5406__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4114_ _4065_/Y _4117_/B _4114_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_68_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_463 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_614 VGND VPWR sky130_fd_sc_hd__decap_12
X_5094_ _5090_/Y _5093_/X _5109_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_110_262 VGND VPWR sky130_fd_sc_hd__decap_12
X_4045_ _4044_/Y _4034_/X _3998_/X _4045_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_56_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4989__A1 _4985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_809 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_883 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3018__A2_N _3017_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5556__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_382 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_842 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4354__A _4340_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_208 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5169__B _5169_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_780 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_599 VGND VPWR sky130_fd_sc_hd__fill_1
X_4947_ _4943_/Y _4946_/X _4947_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_38 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_4878_ _4863_/X _4868_/X _4878_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_166_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_958 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5166__A1 _5165_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3829_ _3829_/A _3806_/X _3829_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_165_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_159 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5185__A _4618_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4913__A1 _4900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_332 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_173 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4529__A _4528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_165 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_809 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3101__B1 _3073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2991__B _2991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_511 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_522 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_382 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_691 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_853 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4264__A _4662_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3476__B1_N _3450_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_730 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_279 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_251 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__A3 _2755_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_441 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_975 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_295 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5157__B2 _5156_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_485 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__A _3608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_479 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_619 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_170 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_97 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_888 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5429__CLK _5429_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_674 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_376 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_739 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_684 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_430 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4439__A _4438_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_964 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3343__A _5470_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_986 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_945 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3062__B _3061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_113 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5579__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_593 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_530 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5093__B1 _5568_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_606 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3997__B _3950_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_691 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4174__A _4172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_886 VGND VPWR sky130_fd_sc_hd__fill_2
X_4801_ _4656_/X _4857_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_739 VGND VPWR sky130_fd_sc_hd__decap_3
X_2993_ _3065_/A _2991_/X _2993_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_21_216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_925 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4902__A _4885_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_62 VGND VPWR sky130_fd_sc_hd__decap_12
X_4732_ _4731_/X _4725_/X data_out2[27] _4726_/X _4732_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_148_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_115 VGND VPWR sky130_fd_sc_hd__fill_2
X_4663_ _4518_/X _4521_/A _4523_/A _4586_/B _3584_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_30_794 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_159 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_3614_ data_in1[2] _3581_/X _3599_/X _3613_/X _3614_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_116_800 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_980 VGND VPWR sky130_fd_sc_hd__fill_2
X_4594_ _5440_/Q _4590_/X _4595_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_116_811 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_822 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2906__B1 _2905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_310 VGND VPWR sky130_fd_sc_hd__fill_1
X_3545_ _2696_/A _3545_/B _3545_/C _3545_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_116_844 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5232__A1_N _5199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_3476_ _5116_/A _3447_/X _3450_/X _3477_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XANTENNA__4659__B1 _4658_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4946__A2_N _4945_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_538 VGND VPWR sky130_fd_sc_hd__decap_8
X_5215_ _5198_/X _5226_/B _5198_/X _5226_/B _5215_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5320__A1 data_in2[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_249 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4349__A _4349_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_750 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3253__A _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5146_ _5143_/X _5145_/Y _5146_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4068__B _4066_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2685__A2 _5366_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_5077_ _5566_/Q _5065_/X _5077_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_319 VGND VPWR sky130_fd_sc_hd__fill_2
X_4028_ _3075_/Y _5537_/Q _3073_/C _3394_/Y _4028_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_25_533 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4084__A _4784_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3398__B1 _4043_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_936 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_232 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_58 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_69 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_939 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_927 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_811 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4250__C _4519_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4898__B1 _4873_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3147__B key_in[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_448 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_855 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_983 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_460 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_482 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5311__A1 _5306_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4259__A _4809_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_709 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3163__A _3028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_62 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_676 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_772 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_219 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3873__A1 _3870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_593 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2796__A2_N _2795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_146 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5093__A2_N _5092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5075__B1 _4942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_937 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_83 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_864 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_897 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_547 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3928__A2 _3837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4722__A _5534_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1014 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_413 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_721 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_231 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_608 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_619 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5544__RESET_B _4309_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_438 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3057__B _3057_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_769 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_3330_ _3254_/Y _3328_/Y _3304_/B _3329_/Y _3330_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_124_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2896__B _2895_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_836 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_3261_ _3291_/A key_in[54] _3261_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4105__A2 _4103_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4169__A _4151_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3073__A _3026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_750 VGND VPWR sky130_fd_sc_hd__fill_2
X_5000_ _5000_/A _4999_/X _5001_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_22_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3192_ _3145_/X key_in[116] _3044_/X _3192_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_79_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_967 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_989 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3801__A _3801_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_499 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_801 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5369__A1 _5300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4632__A _4798_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_878 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3919__A2 _3917_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2976_ _4943_/A _2936_/X _2976_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_147_221 VGND VPWR sky130_fd_sc_hd__decap_12
X_4715_ _5530_/Q _3143_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4592__A2 _4588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3248__A _3201_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_714 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_725 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2874__A1_N _3801_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4646_ _4646_/A _4646_/B _5446_/Q _4645_/X _4646_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_162_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_4577_ _4577_/A _4576_/X _5172_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_3528_ _3528_/A key_in[62] _3528_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_103_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_644 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4079__A _4077_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3459_ _3459_/A _3459_/B _3460_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3414__C _3346_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_379 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5129_ _5129_/A _5129_/B _5130_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3711__A _2717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_477 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_948 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3607__B2 _3606_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3430__B _3431_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_970 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3083__A2 _3057_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2830__A2 _2824_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_333 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4542__A _4542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_700 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_867 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5357__B _5347_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4261__B _4522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_243 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3158__A _3158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_585 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2997__A _2986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_757 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_83 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2897__A2 _2895_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5092__B _5091_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_290 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5523__D _5523_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_952 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_528 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_422 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3846__B2 _3845_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_466 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_989 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5048__B1 _5036_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3621__A _5253_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_285 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_959 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3340__B _3340_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_756 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_458 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_650 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_683 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2821__A2 _2799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_322 VGND VPWR sky130_fd_sc_hd__decap_6
X_2830_ _4637_/X _2824_/X _2825_/X _2826_/X _2829_/X _2830_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__4452__A _4449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5220__B1 _5197_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_221 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5267__B key_in[67] VGND VPWR sky130_fd_sc_hd__diode_2
X_2761_ _2761_/A _2761_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4171__B _4170_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3068__A _3021_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_254 VGND VPWR sky130_fd_sc_hd__fill_2
X_4500_ _4501_/A _4500_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5480_ _3598_/X _5480_/Q _4386_/X _5372_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_416 VGND VPWR sky130_fd_sc_hd__decap_8
X_2692_ _5356_/C _2691_/X _5356_/C _2691_/X _2695_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4431_ _4426_/X _4431_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_717 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5283__A _5252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2700__A _5518_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4362_ _4397_/A _4367_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_300 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_920 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_633 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3515__B _3516_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3313_ _3170_/A _3313_/B _3312_/X _3313_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_99_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_4293_ _4296_/A _4293_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5433__D _4739_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_655 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_3244_ _3244_/A _3244_/B _3244_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3175_ _3175_/A _3175_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4627__A _3337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_477 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_1_0_clock_A clkbuf_4_1_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_447 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3250__B _3249_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_918 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_845 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3557__A1_N _3548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4362__A _4397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4014__A1 _3180_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5466__RESET_B _4402_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_377 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_686 VGND VPWR sky130_fd_sc_hd__decap_12
X_2959_ _2959_/A _3158_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_109_906 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_27 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_522 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_235 VGND VPWR sky130_fd_sc_hd__decap_8
X_4629_ _4518_/X _4629_/B _4578_/A _4629_/D _4630_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_135_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_961 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5193__A _5198_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_588 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3706__A _3704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3525__B1 _3495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_994 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_452 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_42 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_539 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_742 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4537__A _4893_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3441__A _3441_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_285 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4256__B _4658_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_594 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_959 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_296 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_447 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3160__B _3116_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_767 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_650 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_469 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_661 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_806 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3461__C1 _3460_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5368__A _2707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4272__A _4271_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_878 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5202__B1 _5181_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5087__B _5086_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_530 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5518__D _5518_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_563 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_883 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3764__B1 _3748_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_235 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_909 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_543 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3616__A _3606_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_728 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3335__B key_in[56] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_804 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5269__B1 _5267_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_742 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5016__A1_N _5562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_292 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4447__A _4267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_904 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_509 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3295__A2 _3291_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_712 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3070__B _3068_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_756 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_542 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3986__A2_N _3985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_266 VGND VPWR sky130_fd_sc_hd__decap_3
X_4980_ _4968_/X _4971_/X _4980_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_45_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3931_ _3908_/A _3913_/X _3931_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4795__A2 _4674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1001 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_940 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5278__A _5278_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4182__A _4168_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3862_ _3817_/X _3842_/X _3862_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_31_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_675 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_163 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_809 VGND VPWR sky130_fd_sc_hd__decap_3
X_2813_ _2772_/X _2813_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__5428__D _5428_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3793_ _3767_/X _3776_/X _3793_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_118_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_5532_ _5532_/D _3905_/A _4324_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2744_ _5332_/B _5364_/A _2744_/C _2744_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_118_736 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4210__A1_N _4208_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5463_ _5463_/D _5463_/Q _4407_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3526__A _3526_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_599 VGND VPWR sky130_fd_sc_hd__fill_2
X_4414_ _4418_/A _4414_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_172_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_5394_ _4787_/X data_out1[24] _4488_/X _5382_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3245__B _3245_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_653 VGND VPWR sky130_fd_sc_hd__fill_1
X_4345_ _4341_/A _4345_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_59_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_463 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2730__A1 data_in2[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_783 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_314 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_4276_ _4304_/A _4276_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_101_647 VGND VPWR sky130_fd_sc_hd__fill_2
X_3227_ _3227_/A _3226_/X _3227_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4357__A _4354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3481__A1_N _3465_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3261__A _3291_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_168 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3286__A2 _3172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_892 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_3158_ _3158_/A _3158_/B _3159_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_36_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_594 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_380 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_233 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _2889_/Y _3087_/A _3088_/X _3112_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_9 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_620 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4804__B _4803_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_940 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_625 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4092__A _3569_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_973 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_174 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5196__C1 _5195_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_808 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_758 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3436__A _3436_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_52 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_441 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2690__A1_N _5365_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_463 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_260 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2721__B2 _2720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_474 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_923 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5462__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2994__B _2992_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_293 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4267__A reset VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_937 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_469 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5388__RESET_B _4495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_789 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4226__A1 _4225_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_428 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4777__A2 _4769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_748 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_491 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5098__A _5098_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3985__B1 _3957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_995 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_156 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3737__B1 _2771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_863 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3346__A _3343_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_897 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_588 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2960__A1 _2819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2960__B2 _3158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_227 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3065__B _3065_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3504__A3 _3501_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4130_ _4096_/Y _4109_/X _3848_/X _4130_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_69_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_422 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5280__B _5280_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4061_ _4072_/A _4115_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_84_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3268__A2 _3266_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3081__A _5464_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3012_ _3012_/A _3012_/B _3014_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_36_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_767 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_553 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4905__A _4900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_255 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2914__B1_N _2913_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_480 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4768__A2 _4757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_236 VGND VPWR sky130_fd_sc_hd__decap_4
X_4963_ _4870_/X _4961_/Y _4962_/X _2973_/A _4930_/X _5461_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_33_940 VGND VPWR sky130_fd_sc_hd__decap_12
X_3914_ _3909_/X _3912_/Y _3913_/X _3914_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_4894_ _4656_/X _4918_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_634 VGND VPWR sky130_fd_sc_hd__fill_2
X_3845_ _3818_/X _3821_/Y _3817_/X _3845_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_20_678 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4640__A _4639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_511 VGND VPWR sky130_fd_sc_hd__decap_4
X_3776_ _2839_/X _3775_/X _2839_/X _3775_/X _3776_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4997__D _4987_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5515_ _5515_/D _5515_/Q _4344_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_146_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_2727_ _2728_/A _2728_/B _2727_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_146_886 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3256__A _3236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2951__A1 _2989_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5446_ _4613_/Y _5446_/Q _4427_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__5485__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_867 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4153__B1 _4095_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5377_ _4752_/X data_out1[7] _4508_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_472 VGND VPWR sky130_fd_sc_hd__decap_12
X_4328_ _4330_/A _4328_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_86_133 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4087__A _4072_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4259_ _4809_/B _3848_/X _4263_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_74_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_38 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_49 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_789 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4815__A _4815_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4208__A1 _4728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5481__RESET_B _4385_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_87 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5410__RESET_B _4470_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4759__A2 _4757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_98 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_556 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3967__B1 _3966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__C _4519_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_967 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_809 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_617 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4550__A _5553_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2989__B _2989_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3061__B1_N _3060_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_148 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3373__A1_N _3371_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_555 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4931__A2 _4928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_812 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3166__A _3143_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_800 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_834 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_355 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_409 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4695__A1 _2842_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4695__B2 _4688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_899 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_783 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3613__B _3611_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_83 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_764 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5531__D _5531_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5569__RESET_B _4280_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_840 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_756 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_778 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3941__A1_N _3938_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_862 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_169 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4725__A _4699_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_567 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_932 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_792 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_606 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4460__A _4461_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_639 VGND VPWR sky130_fd_sc_hd__fill_2
X_3630_ _3630_/A _3628_/X _3630_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__2899__B key_in[12] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5275__B _5275_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4593__A2_N _4590_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_875 VGND VPWR sky130_fd_sc_hd__fill_2
X_3561_ _3559_/X _3561_/B _3562_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_128_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3076__A _3043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_160 VGND VPWR sky130_fd_sc_hd__fill_1
X_5300_ _5300_/A key_in[36] _5300_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_3492_ data_in2[28] _3391_/X _3462_/X _3491_/Y _5539_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_6_693 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4135__B1 _4133_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5231_ _5481_/Q _5229_/A _5230_/X _5231_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__3804__A _3804_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1005 VGND VPWR sky130_fd_sc_hd__decap_12
X_5162_ _5154_/Y _5156_/X _5160_/B _5169_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__2697__B1 _5356_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4113_ _4068_/A _4113_/B _4117_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_5093_ _5568_/Q _5092_/X _5568_/Q _5092_/X _5093_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__5441__D _4598_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_4044_ _4011_/X _4044_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_84_648 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4989__A2 _4987_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4635__A _4635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_854 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_567 VGND VPWR sky130_fd_sc_hd__decap_12
X_4946_ _4553_/A _4945_/X _4553_/A _4945_/X _4946_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_932 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_606 VGND VPWR sky130_fd_sc_hd__decap_12
X_4877_ _4875_/X _4887_/B _4877_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_166_937 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4370__A _4375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_436 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5166__A2 _5164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3828_ _3828_/A _3805_/Y _3832_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5185__B key_in[64] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_609 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4913__A2 _4899_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3759_ _3759_/A _3758_/X _3759_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_106_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_344 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_558 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_878 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_569 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_141 VGND VPWR sky130_fd_sc_hd__fill_2
X_5429_ _4732_/X data_out2[27] _4446_/X _5429_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_88_910 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_686 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3714__A _3713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_36 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2688__B1 _5343_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_442 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_475 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_64 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3101__A1 data_in2[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_147 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5500__CLK _5429_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_46 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4545__A _4545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_394 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_320 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4264__B _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_191 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_865 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_718 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_23 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_742 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_904 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_56 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_775 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4280__A _4276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_453 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_402 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_947 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_138 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_497 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__B _3607_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_970 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5526__D _3025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_672 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_867 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_355 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_506 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_910 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3624__A _3624_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_837 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_239 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3708__A2_N _3707_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3343__B _3295_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5093__B2 _5092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_467 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4455__A _4469_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3997__C _3010_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_478 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_394 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4174__B _4174_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4800_ _4799_/Y _4800_/B _4813_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_61_353 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2979__A2_N _2978_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_2992_ _3065_/A _2991_/X _2992_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_21_228 VGND VPWR sky130_fd_sc_hd__decap_8
X_4731_ _5538_/Q _4731_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4902__B _4889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5286__A _5256_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_751 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2703__A _5358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_4662_ _4525_/X _4586_/B _4519_/X _4649_/X _4662_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_163_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_3613_ _3579_/A _3611_/X _3612_/Y _3613_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4593_ _5440_/Q _4590_/X _5440_/Q _4590_/X _4593_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__5436__D _4532_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_683 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2906__A1 _4642_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3544_ _3543_/A _3543_/B _3545_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_171_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_631 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_653 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4108__B1 _4107_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_707 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2917__A2_N _2916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_729 VGND VPWR sky130_fd_sc_hd__decap_3
X_3475_ _5128_/A _3474_/X _5128_/A _3474_/X _3475_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5214__A2_N _5213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4659__A1 _4576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_697 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_314 VGND VPWR sky130_fd_sc_hd__decap_12
X_5214_ _5202_/X _5213_/X _5202_/X _5213_/X _5226_/B VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__5320__A2 _5222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3253__B _3253_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5523__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_5145_ _4572_/A _5144_/X _4572_/A _5144_/X _5145_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_57_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_250 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_550 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_475 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_924 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_626 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_572 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2685__A3 _5367_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5076_ _5076_/A _5076_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_57_659 VGND VPWR sky130_fd_sc_hd__fill_2
X_4027_ _4013_/Y _4027_/B _4039_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4365__A _4367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_350 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_501 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4831__A1 _4830_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_843 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_545 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4084__B _4083_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_876 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3398__A1 _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3398__B2 _3397_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4929_ _4928_/A _4927_/X _4929_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_40_559 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_740 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_55 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_948 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_906 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4898__A1 _4908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_20 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_992 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4250__D _4525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_35 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_86 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_472 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_837 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3444__A _3501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5311__A2 _5308_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_633 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_30 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4259__B _3848_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3163__B _3163_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_615 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_85 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3873__A2 _3869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_434 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_294 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5075__A1 _5470_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_862 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_916 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4275__A _4269_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3086__B1 _3875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_670 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_949 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4822__A1 _4821_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2833__B1 _2858_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_876 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_375 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_397 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_403 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3619__A _3619_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_425 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_250 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_745 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_756 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_244 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_778 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_755 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_243 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_788 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_265 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3057__C _3055_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_962 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3017__A2_N _3016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_504 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5546__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3354__A _3354_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3260_ _3259_/A _3258_/Y _3305_/B _3273_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__5513__RESET_B _4346_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_347 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3073__B _2884_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_902 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_369 VGND VPWR sky130_fd_sc_hd__decap_12
X_3191_ _3148_/A key_in[84] _3191_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_78_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_773 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_924 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_103 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_732 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_434 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_1_0_clock_A clkbuf_2_0_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3801__B _3820_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4185__A _4126_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_810 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_821 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_813 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_684 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5369__A2 key_in[102] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2841__A2_N _2840_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2975_ _2913_/A _2938_/X _2975_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3529__A _3529_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4714_ _5529_/Q _4712_/X data_out2[18] _4713_/X _5420_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_147_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_4645_ _4644_/X _4645_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_107_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_428 VGND VPWR sky130_fd_sc_hd__decap_6
X_4576_ _4575_/X _4576_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_269 VGND VPWR sky130_fd_sc_hd__decap_6
X_3527_ _3526_/A _3526_/B _3526_/X _3527_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_115_141 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_515 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_623 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4079__B _4078_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3458_ _3459_/A _3459_/B _3458_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_131_656 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_166 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_870 VGND VPWR sky130_fd_sc_hd__fill_1
X_3389_ _3317_/X _3389_/B _3388_/X _3389_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_97_592 VGND VPWR sky130_fd_sc_hd__decap_6
X_5128_ _5128_/A _5132_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_69_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_147 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_905 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3711__B _3710_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4095__A _4094_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5059_ _5059_/A _5058_/X _5072_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_57_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_692 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_651 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_876 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_353 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4823__A _4823_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_824 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5419__CLK _5413_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_301 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_386 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2830__A3 _2825_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_537 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_98 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4542__B _4542_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_345 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_570 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3240__B1 _3249_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4261__C _4615_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_255 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3158__B _3158_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_575 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5569__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_737 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2997__B _2992_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_258 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_257 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4740__B1 data_out1[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_995 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_51 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_697 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3174__A _3216_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_924 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3902__A _3839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_188 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_592 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_71 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5048__A1 _4896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3621__B _2734_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5048__B2 _4806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3059__B1 _3039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_843 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_982 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_695 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2821__A3 _2752_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5220__A1 data_in2[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3349__A _3349_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2760_ _2759_/X _2761_/A VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2949__A1_N _2998_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_233 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3068__B _3064_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_552 VGND VPWR sky130_fd_sc_hd__decap_12
X_2691_ _5358_/Y _2690_/Y _5358_/Y _2690_/Y _2691_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_299 VGND VPWR sky130_fd_sc_hd__fill_2
X_4430_ _4426_/X _4430_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_759 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5283__B _5252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3534__A1 _5143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_802 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_729 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_770 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_461 VGND VPWR sky130_fd_sc_hd__fill_2
X_4361_ _4267_/Y _4397_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_420 VGND VPWR sky130_fd_sc_hd__decap_12
X_3312_ _3312_/A _3352_/B _3312_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4292_ _4296_/A _4292_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_389 VGND VPWR sky130_fd_sc_hd__decap_8
X_3243_ _3244_/A _3244_/B _3245_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4908__A _4874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3298__B1 _3267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_721 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3812__A _3765_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3174_ _3216_/A _3143_/B _3175_/A _3174_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_66_242 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_787 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_990 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3524__A2_N _3523_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_245 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_5_0_clock_A clkbuf_4_5_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_278 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_993 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_790 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_654 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_317 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4014__A2 _4012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3259__A _3259_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_698 VGND VPWR sky130_fd_sc_hd__decap_4
X_2958_ _3026_/A _2884_/B _2984_/A _2958_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_41_39 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3773__A1 _3769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_2889_ _2889_/A _2889_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_163_534 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_439 VGND VPWR sky130_fd_sc_hd__fill_2
X_4628_ _3501_/A _3529_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5435__RESET_B _4439_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3706__B _3705_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3525__A1 _3178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_973 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3525__B2 _3497_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4559_ _4559_/A _4557_/B _4559_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_1_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_239 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_32 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4818__A _5543_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_54 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_220 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_754 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3441__B _3441_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_873 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_42 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4789__B1 data_out1[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_908 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_673 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4553__A _4553_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3461__B1 _3434_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5368__B key_in[70] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_131 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5391__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3169__A _3169_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5202__B2 _5201_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_890 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_349 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3764__A1 data_in1[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_748 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2801__A _2801_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_940 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_247 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_109 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_984 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3602__A1_N _3588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_781 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5534__D _3314_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_239 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5269__A1 _4636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5269__B2 _5268_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_998 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4728__A _5536_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_916 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3295__A3 _3292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_264 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2873__A1_N _2871_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_554 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_109 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4463__A _4468_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4884__A2_N _4883_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3930_ _3918_/Y _3925_/Y _3945_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_16_172 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5278__B _5278_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_3861_ _3750_/Y _3859_/X _3860_/X _3861_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__4182__B _4182_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_687 VGND VPWR sky130_fd_sc_hd__decap_12
X_2812_ _2733_/A _2698_/B _2842_/A _2812_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_82_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3204__B1 _3217_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_890 VGND VPWR sky130_fd_sc_hd__fill_2
X_3792_ _3681_/A _3794_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_158_873 VGND VPWR sky130_fd_sc_hd__decap_12
X_5531_ _5531_/D _3175_/A _4325_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_2743_ _2719_/A _2718_/A _2743_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_118_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_372 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5294__A _5294_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3807__A _3791_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2711__A _4871_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5462_ _5462_/D _5462_/Q _4408_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4704__B1 data_out2[13] VGND VPWR sky130_fd_sc_hd__diode_2
X_4413_ _4418_/A _4413_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3526__B _3526_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5444__D _5444_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_5393_ _4785_/X data_out1[23] _4489_/X _5498_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_172_397 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_239 VGND VPWR sky130_fd_sc_hd__decap_4
X_4344_ _4341_/A _4344_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_559 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3245__C _3244_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_751 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_976 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_762 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_453 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2730__A2 _5222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_19 VGND VPWR sky130_fd_sc_hd__fill_2
X_4275_ _4269_/A _4304_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_849 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4638__A _4637_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3542__A _3542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_125 VGND VPWR sky130_fd_sc_hd__fill_1
X_3226_ _5468_/Q _3226_/B _3226_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_100_147 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3261__B key_in[54] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_702 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_938 VGND VPWR sky130_fd_sc_hd__fill_1
X_3157_ _3158_/A _3158_/B _3182_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_39_286 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3691__B1 _4750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_448 VGND VPWR sky130_fd_sc_hd__fill_1
X_3088_ _2889_/A _3088_/B _3088_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_716 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_470 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4373__A _4375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_790 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_637 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_687 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_136 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5196__B1 _5175_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_737 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3717__A _3788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_854 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_567 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_943 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_97 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4548__A _4908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_272 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_849 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2994__C _2993_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3452__A _3452_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_307 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_949 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4977__A1_N _4997_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_256 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_565 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4226__A2 _4224_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_50 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4283__A _4304_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_604 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5098__B _5098_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3985__A1 _3958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5529__D _3142_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_687 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5187__B1 _5207_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4934__B1 _4944_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3737__B2 _3736_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_860 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_341 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3346__B _3344_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2960__A2 _2959_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_385 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_613 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4458__A _4461_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3362__A _3317_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_646 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_434 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5111__B1 _5110_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4060_ _4059_/X _4072_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_808 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_145 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_540 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3081__B _3081_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3011_ _2870_/A _3010_/A _3804_/A _3180_/A _3012_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_97_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4193__A2_N _4192_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_757 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_340 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_971 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_727 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3425__B1 _3435_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2706__A _5236_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4962_ _4961_/A _4960_/X _4962_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_952 VGND VPWR sky130_fd_sc_hd__decap_12
X_3913_ _3909_/X _3912_/Y _3913_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__5439__D _4592_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4893_ _4893_/A _5223_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_149_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_136 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4921__A _4873_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3844_ _3842_/X _3843_/Y _3844_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_60_793 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_670 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_3775_ _3773_/X _3774_/X _3775_/X VGND VPWR sky130_fd_sc_hd__xor2_4
X_5514_ _5514_/D _5514_/Q _4345_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2726_ _2726_/A _2728_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_157_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3509__A1_N _3498_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3256__B _3233_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2951__A2 _2989_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5445_ _4612_/X _4646_/B _4428_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_160_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4153__A1 _4073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_879 VGND VPWR sky130_fd_sc_hd__decap_6
X_5376_ _4751_/X data_out1[6] _4509_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_114_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_250 VGND VPWR sky130_fd_sc_hd__fill_2
X_4327_ _4330_/A _4327_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_924 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4368__A _4367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_4258_ _4252_/Y _4615_/B _4258_/C _5576_/D VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_75_819 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_979 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4087__B _4113_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_860 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_478 VGND VPWR sky130_fd_sc_hd__decap_8
X_3209_ _3137_/Y _3209_/B _3209_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_101_489 VGND VPWR sky130_fd_sc_hd__fill_2
X_4189_ _3316_/C _5539_/Q _4188_/X _4189_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_55_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_863 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_407 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4208__A2 _3493_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5199__A _5480_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_930 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3967__A1 _3110_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__D _4253_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_624 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__RESET_B _4422_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_106 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_501 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4550__B _4541_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_512 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_692 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_178 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4931__A3 _4929_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3166__B _3166_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_867 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4695__A2 _4687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4278__A _4276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_581 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3182__A _3160_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3613__C _3612_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_776 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_893 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_381 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3910__A _3860_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_930 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5538__RESET_B _4316_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3958__A1 _3133_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4080__B1 _4050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3308__A2_N _3318_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4741__A _5480_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_478 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_117 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3357__A _3206_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3480__A1_N _3469_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_331 VGND VPWR sky130_fd_sc_hd__fill_2
X_3560_ _3251_/Y _5510_/Q _4791_/X _3397_/Y _3561_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_155_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4239__A1_N _3397_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3076__B key_in[49] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_661 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_684 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_683 VGND VPWR sky130_fd_sc_hd__decap_4
X_3491_ _3317_/X _3491_/B _3490_/X _3491_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_143_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_868 VGND VPWR sky130_fd_sc_hd__fill_2
X_5230_ _3608_/A _2716_/A _5230_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_170_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_193 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4135__B2 _4134_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3804__B _3803_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5161_ _5477_/Q _4995_/X _4542_/B _5160_/X _5477_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4188__A _3980_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_710 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2697__A1 data_in2[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_721 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3894__B1 _3885_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1017 VGND VPWR sky130_fd_sc_hd__decap_3
X_4112_ _4786_/X _4111_/X _4786_/X _4111_/X _4112_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_657 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_5092_ _5052_/A _5091_/X _5092_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4043_ _4026_/A _3950_/B _4043_/C _4043_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_56_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_638 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4916__A _4917_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_830 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3646__B1 _3635_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3820__A _3773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_738 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_866 VGND VPWR sky130_fd_sc_hd__decap_12
X_4945_ _4921_/X _4944_/X _4945_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_52_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_29 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_899 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4651__A _4651_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4876_ _4876_/A _4874_/X _4887_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_21_944 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5452__CLK _5547_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_618 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_977 VGND VPWR sky130_fd_sc_hd__decap_4
X_3827_ _2714_/Y _3825_/X _3826_/Y _3827_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3448__A1_N _5116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3267__A _3344_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_651 VGND VPWR sky130_fd_sc_hd__fill_2
X_3758_ _3756_/X _3757_/X _3756_/X _3757_/X _3758_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_813 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_301 VGND VPWR sky130_fd_sc_hd__decap_4
X_2709_ _4636_/A _2705_/X _2706_/X _2707_/X _2708_/X _2711_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_106_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_621 VGND VPWR sky130_fd_sc_hd__fill_1
X_3689_ _2689_/X _3688_/X _2689_/X _3688_/X _3689_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
X_5428_ _5428_/D data_out2[26] _4449_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_933 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2688__A1 _5335_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5359_ _5490_/Q _2870_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_955 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_465 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_988 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_616 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_329 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3637__B1 _3573_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3730__A _3730_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_297 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_25 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3101__A2 _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_36 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4545__B _4541_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_351 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_811 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_833 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_855 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_332 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4062__B1 _4115_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_376 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_922 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_793 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_410 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4561__A _5562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_398 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_292 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_404 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_465 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_425 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3177__A _4582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_959 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_458 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_835 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_492 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_620 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3905__A _3905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_698 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3624__B _3623_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_890 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5542__D _3567_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3876__B1 _3851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_196 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_605 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_1_0_clock_A clkbuf_2_1_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_830 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4736__A _4699_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5372__RESET_B _4514_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5475__CLK _5574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_2991_ _2988_/X _2991_/B _2991_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_15_782 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4471__A _4475_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4730_ _5537_/Q _4725_/X data_out2[26] _4726_/X _5428_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_159_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_253 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_292 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5286__B _5285_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_106 VGND VPWR sky130_fd_sc_hd__decap_3
X_4661_ _5198_/A _4661_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2703__B _2702_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1010 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3087__A _3087_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3612_ _3609_/X _3610_/Y _3612_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_4592_ _4589_/A _4588_/Y _4591_/Y _4592_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_7_970 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2906__A2 _2903_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3543_ _3543_/A _3543_/B _3545_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_155_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3815__A _3794_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_491 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4108__A1 _4102_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_440 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5305__B1 _5302_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_451 VGND VPWR sky130_fd_sc_hd__decap_6
X_3474_ _4640_/X _3470_/X _3471_/X _3472_/X _3473_/X _3474_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_115_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_827 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4659__A2 _4666_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_518 VGND VPWR sky130_fd_sc_hd__fill_2
X_5213_ _5212_/X _5213_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_495 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5452__D _5452_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_5144_ _5571_/Q _5130_/B _5052_/A _5144_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_69_454 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_638 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4646__A _4646_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5075_ _5470_/Q _4995_/X _4942_/X _5074_/X _5075_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_96_295 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3550__A _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_4026_ _4026_/A _3950_/B _4778_/X _4026_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_37_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4831__A2 _4830_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_833 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_693 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_855 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_696 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3398__A2 _5510_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_398 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4381__A _4381_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4928_ _4928_/A _4927_/X _4928_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_139_916 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_927 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_16 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_735 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_426 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_774 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_89 VGND VPWR sky130_fd_sc_hd__decap_3
X_4859_ _4859_/A _4863_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_138_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_418 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_109 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4898__A2 _4883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_846 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3725__A _3724_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3444__B key_in[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_730 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_645 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_796 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_97 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4556__A _4546_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3460__A _3317_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5498__CLK _5498_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5075__A2 _4995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3086__A1 _2943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3086__B2 _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4822__A2 _4821_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_991 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2833__A1 _4907_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_844 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4035__B1 _3999_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_527 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4291__A _4296_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_562 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_212 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5537__D _5537_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_448 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_256 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_738 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_429 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3546__C1 _3545_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_621 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3057__D _3056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3635__A _3586_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_827 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_461 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3354__B _3309_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3849__B1 _3815_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_337 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3073__C _3073_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3190_ _3148_/A key_in[20] _3190_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_59_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_785 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4466__A _4468_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_744 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_381 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5553__RESET_B _4299_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3370__A _3178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_340 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4185__B _4090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_660 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_395 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_clock_A clkbuf_2_2_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2714__A _2714_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2974_ _2973_/A _2972_/X _2973_/Y _2974_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_148_713 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3529__B key_in[30] VGND VPWR sky130_fd_sc_hd__diode_2
X_4713_ _4701_/A _4713_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5447__D _4807_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_908 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_4644_ _4522_/A _4576_/X _4629_/B _4644_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_162_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_470 VGND VPWR sky130_fd_sc_hd__decap_12
X_4575_ _4518_/X _4524_/Y _4650_/B _4575_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_144_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_492 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3545__A _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3526_ _3526_/A _3526_/B _3526_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_505 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_462 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_409 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_849 VGND VPWR sky130_fd_sc_hd__decap_12
X_3457_ _3488_/A _3457_/B _3459_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_39_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_3388_ _3388_/A _3388_/B _3388_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_112_882 VGND VPWR sky130_fd_sc_hd__decap_3
X_5127_ _4857_/A _5125_/X _5126_/Y _5116_/A _4930_/X _5127_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_58_947 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_733 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4376__A _4397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_958 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_446 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3280__A _4718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_468 VGND VPWR sky130_fd_sc_hd__decap_6
X_5058_ _5030_/Y _5047_/A _5032_/Y _5056_/Y _5057_/X _5058_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_73_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_811 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_38 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4265__B1 all_done VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_822 VGND VPWR sky130_fd_sc_hd__fill_2
X_4009_ _4003_/X _4008_/Y _4009_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_505 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4823__B _4823_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_493 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_357 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5000__A _5000_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_510 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3240__B2 _3239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_704 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_418 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_930 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_237 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3455__A _4731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_974 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4740__A1 _3577_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_665 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4740__B2 _4737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_782 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3174__B _3143_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_933 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3894__A1_N _3885_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_560 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3902__B _3812_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4286__A _4289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_958 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_497 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3190__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_83 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5048__A2 _5046_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_725 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3059__B2 _3058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_693 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_246 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3202__A1_N _3177_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_8 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5220__A2 _4574_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_379 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5513__CLK _5404_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_520 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_908 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_593 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3068__C _3066_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2690_ _5365_/X _2689_/X _5365_/X _2689_/X _2690_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__3847__A1_N _2939_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_92 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_564 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2990__B1 _2950_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_930 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3365__A _3316_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5283__C _5515_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3534__A2 _3504_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4360_ _4354_/X _4360_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_4_12_0_clock_A clkbuf_3_6_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_782 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2742__B1 _2801_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3311_ _3312_/A _3352_/B _3313_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_98_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_101 VGND VPWR sky130_fd_sc_hd__fill_2
X_4291_ _4296_/A _4291_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_140_432 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_3242_ _4718_/X _3280_/B _3241_/X _3244_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3298__A1 _3268_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4908__B _4872_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_178 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3812__B _3812_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_733 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4196__A _4156_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3173_ _5223_/A _3216_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_457 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_928 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4247__B1 _3579_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_696 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_357 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_329 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3259__B _3258_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2957_ _5223_/A _3026_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_4_9_0_clock_A clkbuf_4_9_0_clock/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3773__A2 _3771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_390 VGND VPWR sky130_fd_sc_hd__decap_3
X_2888_ _2999_/A _2887_/X _2888_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_136_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_4627_ _3337_/A _3501_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_163_546 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3275__A _4720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3525__A2 _3495_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4558_ _4987_/A _4557_/B _5560_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_985 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_793 VGND VPWR sky130_fd_sc_hd__decap_3
X_3509_ _3498_/X _3508_/X _3498_/X _3508_/X _3510_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_335 VGND VPWR sky130_fd_sc_hd__decap_4
X_4489_ _4483_/X _4489_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_103_123 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5475__RESET_B _4392_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_476 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5404__RESET_B _4477_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4818__B _4837_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_66 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4238__B1 _4236_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_32 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4789__A1 _4788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4834__A _4833_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4789__B2 _4782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5306__A1_N _4836_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_460 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3016__A2_N _3015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_994 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3461__A1 data_in2[27] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4553__B _4547_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_622 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5536__CLK _5530_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_30 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3646__A2_N _3645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3169__B _3169_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3764__A2 _3697_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_727 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2972__B1 _2970_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_523 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2801__B _2801_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3185__A _3112_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_911 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2724__B1 _2776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_589 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_495 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_966 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3913__A _3909_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5269__A2 _5265_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_733 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5550__D _5550_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_766 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4229__B1 _3523_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_641 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_566 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_780 VGND VPWR sky130_fd_sc_hd__fill_2
X_3860_ _3750_/Y _3859_/X _3860_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_806 VGND VPWR sky130_fd_sc_hd__decap_12
X_2811_ data_in2[9] _2731_/X _2783_/X _2810_/Y _2811_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_60_986 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3204__A1 _3175_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_699 VGND VPWR sky130_fd_sc_hd__decap_3
X_3791_ _3780_/A _3786_/Y _3791_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_31_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_840 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__decap_3
X_5530_ _3171_/X _5530_/Q _4327_/X _5530_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2742_ _5292_/X _2739_/B _2801_/A _2742_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_157_351 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_727 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_513 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3807__B _3806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5294__B _5294_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_395 VGND VPWR sky130_fd_sc_hd__fill_2
X_5461_ _5461_/D _2973_/A _4409_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2711__B _2711_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3095__A _3095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_4412_ _4419_/A _4418_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4704__A1 _2989_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4704__B2 _4701_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5392_ _5392_/D data_out1[22] _4491_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_611 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2715__B1 _5260_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4343_ _4341_/A _4343_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_125_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_508 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5409__CLK _5402_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_251 VGND VPWR sky130_fd_sc_hd__fill_2
X_4274_ _4271_/A _4274_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3542__B _3540_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3225_ _5468_/Q _3226_/B _3227_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__5460__D _4953_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3156_ _3012_/A _3155_/A _3895_/A _3155_/Y _3158_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_55_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_500 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_360 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3691__B2 _3690_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5559__CLK _5555_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4654__A _4525_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3087_ _3087_/A _3088_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_728 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_611 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_482 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_644 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_953 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_806 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_17 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_986 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5196__A1 data_in2[0] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3989_ _3939_/X _3988_/X _3953_/X _3989_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_10_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3717__B _3715_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_332 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_132 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3733__A _3705_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_785 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4548__B _4547_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_284 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_338 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_349 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5370__D _4740_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_42 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_371 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4564__A _5065_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_268 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_942 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3985__A2 _3962_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_666 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_452 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_103 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5187__A1 _5203_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_114 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_137 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_699 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3908__A _3908_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2812__A _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4934__B2 _4933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_872 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_83 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5545__D _4541_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_855 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5397__RESET_B _4485_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3346__C _3345_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_549 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3643__A _3642_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_806 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_828 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_305 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_625 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3362__B _3362_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5111__A1 _5086_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3538__A2_N _3537_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3010_ _3010_/A _3180_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3122__B1 _3120_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4474__A _4475_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_739 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3425__A1 _3395_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2706__B key_in[7] VGND VPWR sky130_fd_sc_hd__diode_2
X_4961_ _4961_/A _4960_/X _4961_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_51_227 VGND VPWR sky130_fd_sc_hd__fill_2
X_3912_ _3889_/Y _3910_/Y _3912_/C _3912_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_33_964 VGND VPWR sky130_fd_sc_hd__decap_12
X_4892_ _4882_/A _4847_/X _4531_/X _4891_/Y _5455_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_32_441 VGND VPWR sky130_fd_sc_hd__fill_2
X_3843_ _3721_/Y _3841_/X _3843_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_149_148 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2722__A _2722_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3774_ _3724_/X _3752_/X _3735_/Y _3636_/Y _3751_/X _3774_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_20_669 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_811 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2936__B1 _2934_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5513_ _5513_/D _5513_/Q _4346_/X _5404_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_9_681 VGND VPWR sky130_fd_sc_hd__decap_12
X_2725_ _5356_/C _2691_/X _2694_/X _2726_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__5455__D _5455_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_803 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_354 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_814 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_5444_ _5444_/D _4646_/A _4429_/X _5469_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4689__B1 data_out2[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4153__A2 _4152_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_5375_ _5375_/D data_out1[5] _4510_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4649__A _4577_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4326_ _4340_/A _4330_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_560 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_582 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_936 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_496 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_947 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5381__CLK _5382_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4257_ _4517_/Y _4667_/X _4256_/X _4258_/C VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_47_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_3208_ _3144_/A _3166_/X _3210_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_28_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_4188_ _3980_/Y _3463_/Y _4188_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4861__B1 _4873_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3139_ _3139_/A _3138_/X _3139_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_55_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_853 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4384__A _4387_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_257 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_363 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_897 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_27 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4613__B1 _5446_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_290 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3967__A2 _3965_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_986 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_958 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_794 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3728__A _3728_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_833 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_855 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5490__RESET_B _4374_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_97 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_869 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4559__A _4559_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3463__A _5539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_614 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_251 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_625 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3182__B _3182_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_113 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_1_1_0_clock_A clkbuf_0_clock/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_511 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3910__B _3888_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4294__A _4296_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_385 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4604__B1 _4603_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_396 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3958__A2 _3956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4080__A1 _4052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_457 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5578__RESET_B _4271_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3638__A _5284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_956 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_619 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_822 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5507__RESET_B _4353_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3357__B _3357_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_844 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3591__B1 _3573_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_505 VGND VPWR sky130_fd_sc_hd__decap_6
X_3490_ _3489_/A _3541_/C _3490_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_155_696 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4469__A _4469_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_912 VGND VPWR sky130_fd_sc_hd__decap_3
X_5160_ _4918_/A _5160_/B _5160_/C _5160_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_151_880 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4188__B _3463_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2697__A2 _5222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_593 VGND VPWR sky130_fd_sc_hd__decap_8
X_4111_ _4096_/Y _4109_/X _4095_/X _4152_/A _4111_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3894__B2 _3893_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_5091_ _4566_/A _5077_/X _5091_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_232 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_989 VGND VPWR sky130_fd_sc_hd__decap_12
X_4042_ data_in1[21] _3976_/X _4026_/X _4041_/Y _4042_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_49_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4916__B _4915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3646__B2 _3645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3820__B _3820_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_842 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2717__A _2717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_190 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_341 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_536 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_193 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4932__A _5554_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_878 VGND VPWR sky130_fd_sc_hd__decap_3
X_4944_ _4944_/A _4932_/X _4944_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_4875_ _4876_/A _4874_/X _4875_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_166_917 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_282 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_591 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3548__A _5542_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_800 VGND VPWR sky130_fd_sc_hd__decap_4
X_3826_ _2714_/Y _3825_/X _3826_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_119_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_3757_ _3587_/B _3737_/X _3720_/Y _3757_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_134_825 VGND VPWR sky130_fd_sc_hd__decap_12
X_2708_ _5299_/A key_in[103] _5303_/A _2708_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_161_611 VGND VPWR sky130_fd_sc_hd__fill_2
X_3688_ _3685_/X _3686_/Y _3687_/X _3688_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_145_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_869 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4379__A _4381_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_5427_ _5427_/D data_out2[25] _4450_/X _5424_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_133_357 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3283__A _3284_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_880 VGND VPWR sky130_fd_sc_hd__fill_1
X_5358_ _5358_/A _5357_/X _5358_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__2688__A2 _2769_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_891 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_593 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_293 VGND VPWR sky130_fd_sc_hd__decap_4
X_4309_ _4305_/A _4309_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_967 VGND VPWR sky130_fd_sc_hd__decap_8
X_5289_ _3578_/A _5288_/A _3577_/A _2799_/A _5290_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_102_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_628 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3637__A1 _5178_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_799 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3637__B2 _3636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_609 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_514 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4842__A _4830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4062__A1 _4043_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_733 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_219 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4561__B _4561_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_766 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3555__A1_N _5164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3458__A _3459_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_788 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_928 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_967 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_276 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_30 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_477 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_85 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3177__B _3176_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_448 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_961 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4192__A2_N _4191_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_471 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4289__A _4289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_654 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3876__A1 _3826_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_422 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3921__A _3873_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_522 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_533 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_341 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_834 VGND VPWR sky130_fd_sc_hd__fill_2
X_2990_ _2930_/A _2989_/X _2950_/X _2991_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_15_761 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_260 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_906 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3368__A _3368_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_276 VGND VPWR sky130_fd_sc_hd__decap_4
X_4660_ _5256_/A _5198_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_30_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_797 VGND VPWR sky130_fd_sc_hd__fill_2
X_3611_ _3609_/X _3610_/Y _3611_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4591_ _4590_/X _4591_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_127_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_994 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_3542_ _3542_/A _3540_/X _3541_/Y _3543_/B VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_116_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4108__A2 _4105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3815__B _3814_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_858 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5305__A1 _4637_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_964 VGND VPWR sky130_fd_sc_hd__decap_12
X_3473_ _3499_/A key_in[124] _3408_/X _3473_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4199__A _4159_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_869 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5305__B2 _5304_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_817 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_154 VGND VPWR sky130_fd_sc_hd__decap_3
X_5212_ _5211_/A _5210_/X _5211_/X _5212_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_115_379 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_731 VGND VPWR sky130_fd_sc_hd__fill_1
X_5143_ _5143_/A _5143_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4927__A _4911_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3831__A _3831_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_786 VGND VPWR sky130_fd_sc_hd__fill_2
X_5074_ _5071_/Y _5072_/X _5073_/Y _5074_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_111_585 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4816__B1 _5448_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4646__B _4646_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_959 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_596 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3550__B key_in[63] VGND VPWR sky130_fd_sc_hd__diode_2
X_4025_ data_in1[20] _3976_/X _3997_/X _4024_/Y _5499_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_37_330 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_801 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_812 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_396 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_709 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4662__A _4525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5429__RESET_B _4446_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4927_ _4911_/X _4917_/X _4927_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_21_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_4858_ _4848_/A _4847_/X _4531_/X _4857_/X _5452_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_60_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_747 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_438 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_3809_ _3788_/A _3807_/Y _3808_/X _3809_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_4789_ _4788_/X _4781_/X data_out1[25] _4782_/X _5395_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_107_803 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_407 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3555__B1 _5164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2910__A _2907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_324 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_953 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_452 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_986 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_463 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3307__B1 _3299_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_602 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_230 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4837__A _5543_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_861 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3307__A2_N _3306_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4223__A1_N _3395_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3741__A _3741_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_105 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_959 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4807__B1 _4798_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_831 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3460__B _3458_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3086__A2 _4043_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_160 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2833__A2 _2830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_631 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_193 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4572__A _4572_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4035__A1 _3848_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5232__B1 _5181_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_686 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_539 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_185 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_574 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_764 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_775 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_769 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_274 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_268 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3916__A _3904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3546__B1 _3519_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_920 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_482 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3635__B _3634_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5553__D _5553_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_463 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_305 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_880 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3849__A1 _3848_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1004 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3651__A _3651_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5442__CLK _5469_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_959 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3370__B _3369_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4185__C _3300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_992 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_642 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4482__A _4477_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_973 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5522__RESET_B _4336_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_528 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_2973_ _2973_/A _2972_/X _2973_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_148_703 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3098__A _3099_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4712_ _4699_/A _4712_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4643_ _4616_/X _4641_/X _4642_/Y _4616_/X _4643_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_163_706 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_717 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_268 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3826__A _2714_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3537__B1 _3522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_983 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_4574_ _5165_/A _4574_/B _4574_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_128_482 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1010 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3545__B _3545_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3525_ _3178_/Y _3495_/B _3495_/X _3497_/X _3526_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__5463__D _5463_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_666 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_986 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_603 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_474 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_3456_ _4731_/X _3455_/B _3457_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_131_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4657__A _4629_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3387_ _3388_/A _3388_/B _3389_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_97_550 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3561__A _3559_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5271__B1_N _5270_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_5126_ _5125_/A _5124_/X _5126_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_57_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_745 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3280__B _3280_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_5057_ _5028_/Y _5057_/B _5057_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4265__A1 _4629_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_108 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_992 VGND VPWR sky130_fd_sc_hd__decap_12
X_4008_ _3983_/Y _4008_/B _4006_/Y _4007_/Y _4008_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_72_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_940 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4392__A _4390_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2905__A _2905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5214__B1 _5202_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_517 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_483 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_848 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_859 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5000__B _4999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3776__B1 _2839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_544 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_235 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_909 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_216 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_920 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_953 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3455__B _3455_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4740__A2 _4736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5373__D _5373_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_474 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_614 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5465__CLK _5579_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3174__C _3175_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_198 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4567__A _5568_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_977 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3471__A _3501_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_872 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3902__C _3902_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_691 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3190__B key_in[20] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5048__A3 _5047_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_95 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4177__A1_N _4171_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_737 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_480 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_642 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2815__A _5358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_837 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5548__D _5548_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_500 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_202 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_213 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_544 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3068__D _3067_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2990__A1 _2930_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_249 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3365__B _3365_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4192__B1 _3479_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_760 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2742__A1 _5292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_923 VGND VPWR sky130_fd_sc_hd__fill_2
X_3310_ _3287_/C _3309_/B _3309_/Y _3352_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_153_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_271 VGND VPWR sky130_fd_sc_hd__decap_4
X_4290_ _4304_/A _4296_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_152_293 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_281 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_124 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_292 VGND VPWR sky130_fd_sc_hd__decap_4
X_3241_ _4718_/X _3280_/B _3241_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4477__A _4477_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3298__A2 _3271_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4908__C _4908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_572 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3812__C _2714_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3172_ _5222_/A _3172_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4196__B _4196_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_778 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4247__A1 _4246_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_715 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_597 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_631 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_826 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5101__A _5568_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_303 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_494 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5458__D _5458_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_859 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3758__B1 _3756_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_369 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4940__A _4918_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2956_ _5222_/A _2956_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_544 VGND VPWR sky130_fd_sc_hd__decap_4
X_2887_ _2887_/A _2887_/B _2887_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3556__A _3556_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_739 VGND VPWR sky130_fd_sc_hd__decap_12
X_4626_ _3293_/A _3337_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__5488__CLK _5372_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3275__B _3274_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_430 VGND VPWR sky130_fd_sc_hd__decap_12
X_4557_ _4997_/C _4557_/B _5559_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_463 VGND VPWR sky130_fd_sc_hd__fill_2
X_3508_ _3505_/X _3507_/B _3507_/X _3508_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_143_271 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_282 VGND VPWR sky130_fd_sc_hd__decap_4
X_4488_ _4483_/X _4488_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_23 VGND VPWR sky130_fd_sc_hd__decap_8
X_3439_ _4784_/X _4791_/X _3108_/A _3251_/A _3441_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4387__A _4387_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3291__A _3291_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_89 VGND VPWR sky130_fd_sc_hd__decap_3
X_5109_ _5082_/Y _5109_/B _5109_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4238__A1 _3523_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5444__RESET_B _4429_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_970 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_886 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_586 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_620 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_439 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4834__B _4833_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4789__A2 _4781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_804 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_152 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5011__A _4891_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3461__A2 _3391_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_809 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_667 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4850__A _4819_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_318 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_352 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3466__A _3155_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2972__A1 _4637_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2972__B2 _2971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_385 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_920 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3185__B _3185_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_579 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2724__A1 _2723_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_997 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_934 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_945 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3913__B _3912_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_741 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5269__A3 _5266_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4297__A _4304_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_723 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_73 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_273 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_778 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_789 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4229__B2 _4228_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_409 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_664 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_995 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_792 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_185 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_133 VGND VPWR sky130_fd_sc_hd__fill_2
X_2810_ _2852_/A _2808_/Y _2809_/X _2810_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_20_818 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4760__A _5490_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3790_ _3765_/A _3679_/B _3804_/A _3790_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3204__A2 _3203_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_881 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_852 VGND VPWR sky130_fd_sc_hd__fill_2
X_2741_ _2741_/A _2801_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_158_886 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3376__A _3337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_525 VGND VPWR sky130_fd_sc_hd__decap_3
X_5460_ _4953_/X _4943_/A _4410_/X _5555_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_68_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_709 VGND VPWR sky130_fd_sc_hd__decap_4
X_4411_ _4411_/A _4411_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4704__A2 _4699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_366 VGND VPWR sky130_fd_sc_hd__decap_6
X_5391_ _4779_/X data_out1[21] _4492_/X _5574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2715__A1 _3626_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2715__B2 _2714_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_4342_ _4341_/A _4342_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_28_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_656 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_4273_ _4271_/A _4273_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_466 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_200 VGND VPWR sky130_fd_sc_hd__decap_4
X_3224_ _4638_/X _3218_/X _3219_/X _3220_/X _3223_/X _3226_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__3542__C _3541_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4000__A _5536_/Q VGND VPWR sky130_fd_sc_hd__diode_2
.ends


* NGSPICE file created from usb.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 D Q RESET_B CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 D Q SET_B CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 D Q CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

.subckt usb clk_48 data_in[0] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5]
+ data_in[6] data_in[7] data_in_valid data_out[0] data_out[1] data_out[2] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] data_strobe data_toggle direction_in
+ endpoint[0] endpoint[1] endpoint[2] endpoint[3] handshake[0] handshake[1] rst_n
+ rx_j rx_se0 setup success transaction_active tx_en tx_j tx_se0 usb_address[0] usb_address[1]
+ usb_address[2] usb_address[3] usb_address[4] usb_address[5] usb_address[6] usb_rst
+ VPWR VGND
XFILLER_39_222 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1151__B1 _1158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_133 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1206__B2 _1205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1206__A1 _1214_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0965__B1 _1447_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1390__B1 _1389_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__D handshake[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1147__C _1147_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1270_ _1363_/A _1247_/D _1270_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_70 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1133__B1 _1147_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_217 VGND VPWR sky130_fd_sc_hd__fill_2
X_0985_ _0979_/X _0980_/X _1444_/Q data_out[1] _0981_/X _0985_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_8_170 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1004__A1_N _1552_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1606_ _1417_/Y _1606_/Q rst_n _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_1537_ _1537_/D _1537_/Q _0927_/X _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1372__B1 _0769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1354__A data_in_valid VGND VPWR sky130_fd_sc_hd__diode_2
X_1468_ _1467_/Q _0766_/A _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1504__D _1504_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1399_ data_in[6] _1399_/B _1399_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_27_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1248__B _1245_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_280 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_50 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_272 VGND VPWR sky130_fd_sc_hd__fill_2
X_0770_ _0716_/X _0887_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1158__B _1155_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0997__B _0816_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_125 VGND VPWR sky130_fd_sc_hd__fill_2
X_1322_ _0869_/A _1358_/A _1322_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1253_ _1241_/X _1251_/Y _1252_/X _1607_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_64_353 VGND VPWR sky130_fd_sc_hd__decap_3
X_1184_ _1095_/X _1183_/X _1181_/X _1184_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_24_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0865__C1 _0864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_250 VGND VPWR sky130_fd_sc_hd__fill_2
X_0968_ _0855_/X _0955_/X _1442_/Q _1450_/Q _0958_/X _0968_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_0899_ _1358_/A _0892_/X _0894_/X _0898_/X _0899_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1345__B1 _1330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1084__A _1550_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_239 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1250__C _1250_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_53 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1259__A _1250_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_334 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0735__A1_N usb_address[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_261 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1442__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0822_ _0821_/Y _0823_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0753_ _0734_/Y _0753_/B _0742_/X _0753_/D _0754_/D VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0801__A _0799_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1592__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1569__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_1305_ _1305_/A _1305_/B _0712_/B _1306_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_37_331 VGND VPWR sky130_fd_sc_hd__fill_2
X_1236_ _1603_/Q _1236_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_1167_ _0916_/A _1160_/X _1167_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_397 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_1098_ _1555_/Q _1094_/X _1556_/Q _1095_/X _1098_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_52_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0711__A _1305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1030__A2 _0853_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1097__A2 _1094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1465__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_356 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_367 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1536__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_389 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1599__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1088__A2 _1059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1021_ _0998_/X _1021_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_19_375 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1602__D _1235_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_397 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_389 VGND VPWR sky130_fd_sc_hd__fill_2
X_0805_ _1466_/Q _1466_/D _0798_/A _0805_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0736_ _1529_/Q _0736_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_29_117 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1362__A _0715_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1512__D _1512_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1219_ _1200_/A _1222_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_55_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1079__A2 _1069_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_150 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1488__CLK _1514_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_334 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_161 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1279__A2_N _1278_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0706__A _0759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1251__A2 _1244_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1272__A _1272_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_183 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1422__D _1422_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_6_0_clk_48_A clkbuf_4_7_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_378 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_175 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_359 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_23 VGND VPWR sky130_fd_sc_hd__fill_2
X_1570_ _1570_/D _0918_/B rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_6_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_260 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1182__A _1183_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1004_ _1552_/Q _0840_/X _1552_/Q _0840_/X _1004_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1584__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1233__A2 _1205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1513__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__C _0894_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1357__A _1350_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1076__B _1064_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1507__D _1507_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0719_ _0719_/A _0718_/X _0719_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_223 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1092__A _1095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_278 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_142 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_123 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1503__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_381 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0983__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0983__B2 _0981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1267__A _1272_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__B2 _1447_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_230 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_223 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_237 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1215__A2 _1208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_178 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1281__A1_N _1272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0974__A1 _0969_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0974__B2 _0972_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_1553_ _1553_/D _0904_/A rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1484_ _1484_/D _1484_/Q rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1151__A1 _1149_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_278 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1526__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_167 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1206__A2 _1204_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0965__B2 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0965__A1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_clk_48_A clkbuf_3_6_0_clk_48/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1390__A1 _1388_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_79 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1133__A1 _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1549__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1610__D _1303_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_229 VGND VPWR sky130_fd_sc_hd__decap_3
X_0984_ _0979_/X _0980_/X _1443_/Q data_out[0] _0981_/X _1427_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_8_193 VGND VPWR sky130_fd_sc_hd__fill_2
X_1605_ _1605_/D _1605_/Q rst_n _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1536_ _1054_/X _1536_/Q _0927_/X _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1372__A1 _1409_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1354__B _0887_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1467_ rx_j _1467_/Q _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1124__A1 _1566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1398_ _0887_/A _0758_/Y data_in[5] _1424_/Q _1397_/X _1424_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1370__A _1369_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1520__D _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0714__A _0714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_11 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_148 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1060__B1 _1056_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1248__C _0874_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1115__A1 _0919_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1430__D _1430_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_73 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1158__C _1158_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0997__C _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1605__D _1605_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1321_ _0780_/A _0795_/X _1321_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_1_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_1252_ _1252_/A _1252_/B _1252_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_64_321 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1190__A _0717_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1183_ _1587_/Q _1183_/B _1183_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_49_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0865__B1 _1319_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_284 VGND VPWR sky130_fd_sc_hd__decap_3
X_0967_ _0747_/Y _0962_/Y _1441_/Q _0962_/Y _0967_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1042__B1 _0825_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0898_ _1492_/Q _0898_/B _0898_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1365__A _0869_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1345__A1 _0772_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1084__B _1014_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1519_ _1519_/D _0755_/B rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1515__D _1328_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_192 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0709__A _1606_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_218 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_229 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1250__D _1254_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1281__B1 _0707_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1259__B _0874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1033__B1 _0755_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1425__D _1425_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_72 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_357 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_34 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_89 VGND VPWR sky130_fd_sc_hd__decap_4
X_0821_ _0994_/A _0821_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1024__B1 _1522_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0752_ _0744_/X _0746_/X _0749_/X _0751_/Y _0753_/D VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0801__B _0800_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1185__A _1470_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1304_ _1305_/A _1296_/X _0712_/B _1304_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_56_107 VGND VPWR sky130_fd_sc_hd__fill_2
X_1235_ _1601_/Q _1205_/X _1234_/X _1235_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_49_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_1166_ _1165_/X _1166_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0842__A1_N _0837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_376 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_173 VGND VPWR sky130_fd_sc_hd__decap_4
X_1097_ _1554_/Q _1094_/X _1555_/Q _1095_/X _1097_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1263__B1 _1250_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1015__B1 _1529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1095__A _1095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_321 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_398 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_20 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_64 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_86 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_236 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0902__A _0810_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_107 VGND VPWR sky130_fd_sc_hd__fill_2
X_1020_ _0823_/B _1020_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_19_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_368 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_195 VGND VPWR sky130_fd_sc_hd__decap_4
X_0804_ _0797_/Y _0802_/X _0803_/X _0808_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0812__A _1583_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_280 VGND VPWR sky130_fd_sc_hd__fill_2
X_0735_ usb_address[4] _1447_/Q usb_address[4] _1447_/Q _0753_/B VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__1542__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1362__B _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_1218_ _1593_/Q _1216_/X _1217_/X _1218_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_37_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_1149_ _1148_/Y _1149_/B _1149_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_37_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_305 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_206 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0722__A _0721_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0734__A1_N usb_address[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1432__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_162 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1582__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1227__B1 _1226_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_327 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_272 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1163__C1 _1162_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_235 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1182__B _1181_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1003_ _1003_/A _1086_/A _1550_/Q _1003_/D _1005_/C VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_19_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1218__B1 _1217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__D _0898_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1357__B _1357_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0718_ _0717_/X _0718_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1553__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1455__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1373__A _0725_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1523__D _1523_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0717__A _0717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1209__B1 _1589_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_371 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0983__A2 _0980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1393__C1 _1392_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1433__D _0990_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_320 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0974__A2 _0971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1478__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1608__D _1257_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1552_ _1552_/D _1552_/Q _0927_/X _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1483_ _1312_/X _1309_/A _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1193__A _0873_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1151__A2 _1150_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_308 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_319 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0965__A2 _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1518__D _1518_/D VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0_clk_48 clkbuf_0_clk_48/X clkbuf_2_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1390__A2 _1362_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_64 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1428__D _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0910__A _0909_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1133__A2 _1130_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0983_ _0979_/X _0980_/X _1527_/Q _1442_/Q _0981_/X _0983_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__0820__A _1102_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1604_ _1239_/X _1604_/Q _0928_/X _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1535_ _1053_/X _1013_/C _0927_/X _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1372__A2 _0889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1354__C _0757_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1466_ _1466_/D _1466_/Q _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1124__A2 _1120_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1397_ _1364_/X _1397_/B _1397_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_27_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_252 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_138 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1060__A1 _1056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1060__B2 _1004_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_304 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0730__A _1317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1348__C1 _1330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_341 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1115__A2 _1111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_97 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0905__A _1556_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_131 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_164 VGND VPWR sky130_fd_sc_hd__fill_2
X_1320_ _1315_/Y _0794_/Y _1319_/X _0870_/Y _1504_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__1516__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1251_ _1252_/A _1244_/X _1247_/X _1248_/X _1250_/X _1251_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
X_1182_ _1183_/B _1181_/X _1182_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__0865__A1 _1492_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1190__B _1186_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_219 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0815__A _0810_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0966_ _0855_/X _0955_/X _1440_/Q _0744_/B _0958_/X _0966_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1042__B2 _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1042__A1 _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0897_ _1316_/B _0895_/X _0732_/A _0896_/X _0898_/B VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__1365__B _0872_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_19 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1345__A2 _1339_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_127 VGND VPWR sky130_fd_sc_hd__fill_1
X_1518_ _1518_/D _1317_/A rst_n _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1449_ _0967_/X _1449_/Q _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_4_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_300 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1381__A _1381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_333 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0709__B _1605_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1531__D _0995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0725__A _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1281__B2 _1240_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_33 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1033__B2 _0853_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1033__A1 _0837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1539__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1047__A2_N _1010_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_333 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1441__D _0982_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0847__A1 _1485_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_377 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_clk_48 clkbuf_2_3_0_clk_48/A clkbuf_3_7_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1490__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_296 VGND VPWR sky130_fd_sc_hd__fill_2
X_0820_ _1102_/A _1187_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1024__A1 _1020_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1024__B2 _1021_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0751_ _0745_/Y _1444_/Q _0750_/X _0751_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1185__B _1185_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clk_48_A clkbuf_2_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1303_ _1303_/A _1298_/X _1302_/Y _1303_/X VGND VPWR sky130_fd_sc_hd__and3_4
Xclkbuf_4_11_0_clk_48 clkbuf_3_5_0_clk_48/X _1609_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1234_ _1234_/A _1200_/A _1234_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1165_ _1164_/X _1165_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1578__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_1096_ _0904_/A _1094_/X _1554_/Q _1095_/X _1554_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1507__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk_48 clk_48 clkbuf_0_clk_48/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_20_200 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1263__A1 _1252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_288 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1015__A1 _1533_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1015__B2 _0996_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0949_ endpoint[1] _0945_/B _0949_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1526__D _1028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_355 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0964__A1_N _0740_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_54 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_200 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_97 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1436__D _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_163 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_199 VGND VPWR sky130_fd_sc_hd__fill_2
X_0803_ _0799_/Y _0800_/Y _0798_/Y _0802_/B _0803_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1196__A _1196_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0734_ usb_address[0] _1443_/Q usb_address[0] _1443_/Q _0734_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_6_292 VGND VPWR sky130_fd_sc_hd__fill_2
X_1217_ _1217_/A _1214_/B _1217_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_25_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_1148_ _1573_/Q _1148_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_25_358 VGND VPWR sky130_fd_sc_hd__fill_2
X_1079_ _1002_/C _1069_/X _1078_/X _1079_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_40_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0995__B1 _0993_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_21 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1227__A1 _1597_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0986__B1 data_out[2] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1163__B1 _1147_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_258 VGND VPWR sky130_fd_sc_hd__fill_2
X_1002_ _1072_/A _1078_/A _1002_/C _1002_/D _1003_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_19_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_144 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1218__A1 _1593_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0823__A _0823_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0977__B1 _1439_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_394 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1357__C _1329_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0717_ _0717_/A _1470_/Q _0717_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1373__B _1372_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_clk_48 clkbuf_3_7_0_clk_48/A clkbuf_3_6_0_clk_48/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_57_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1522__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0717__B _1470_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1209__B2 _1208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0733__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0968__B1 _1450_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0983__A3 _1527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1393__B1 _1386_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0908__A _1557_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_122 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_114 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_361 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0959__B1 _1443_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0974__A3 _1521_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_1551_ _1551_/D _1086_/A _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1482_ _1293_/Y _1482_/Q _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_39_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_206 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0818__A _1102_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1422__CLK _1514_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0965__A3 _1439_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1384__A data_in[2] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1572__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1534__D _1052_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0728__A _0777_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_280 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_272 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1366__B1 _1410_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_309 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1444__D _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_51 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1445__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0982_ _0979_/X _0980_/X _1526_/Q _1441_/Q _0981_/X _0982_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_8_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1595__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1603_ _1237_/X _1603_/Q _0928_/X _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1534_ _1052_/Y _1534_/Q _0927_/X _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1465_ _0806_/A _1466_/D _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1396_ _1423_/Q _1394_/X _1373_/Y _1395_/X _1396_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_35_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1379__A _1315_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1529__D _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1060__A2 _1059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1348__B1 _1347_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0730__B _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_32 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_228 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_239 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1468__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_250 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_clk_48_A clkbuf_3_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1277__A2_N _1276_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1289__A _1406_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_253 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_97 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_clk_48 clkbuf_4_9_0_clk_48/A _1514_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_41_297 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1439__D _1439_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0921__A _1567_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_176 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_7 VGND VPWR sky130_fd_sc_hd__fill_1
X_1250_ _1250_/A _1245_/X _1250_/C _1254_/D _1250_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_49_331 VGND VPWR sky130_fd_sc_hd__fill_1
X_1181_ _1588_/Q _1187_/B _1181_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_49_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0865__A2 _0879_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_261 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0815__B _0909_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1199__A _1205_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0965_ _0855_/X _0955_/X _1439_/Q _1447_/Q _0958_/X _1447_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1042__A2 _0837_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0896_ _1313_/A _0794_/B _0776_/B _0896_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_1517_ _1031_/X _0776_/B rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1448_ _0966_/X _0744_/B _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1610__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1381__B _0722_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1379_ _1315_/A _0786_/Y _1380_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_367 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0725__B _0725_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1033__A2 _0853_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_179 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_183 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0847__A2 _0818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_315 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0916__A _0916_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_389 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__A2 _0825_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0750_ usb_address[2] _0738_/Y _0750_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_1302_ _1301_/X _1302_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_1233_ _1600_/Q _1205_/X _1232_/X _1233_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_29_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_172 VGND VPWR sky130_fd_sc_hd__decap_3
X_1164_ _0916_/A _1160_/X _1164_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_37_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0826__A _0994_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1095_ _1095_/A _1095_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_52_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1263__A2 _1262_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_234 VGND VPWR sky130_fd_sc_hd__decap_4
X_0948_ _1450_/Q _0942_/X _0947_/X _1497_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1015__A2 _1010_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0879_ _0879_/A _0879_/B _0879_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__1392__A _0886_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1542__D _1068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_142 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_345 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0736__A _1529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_389 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1506__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_43 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_85 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1452__D _1415_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_304 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_392 VGND VPWR sky130_fd_sc_hd__decap_4
X_0802_ _0798_/Y _0802_/B _0802_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0733_ _0733_/A _0862_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1216_ _1205_/A _1216_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_37_142 VGND VPWR sky130_fd_sc_hd__fill_2
X_1147_ _1147_/A _1149_/B _1147_/C _1572_/D VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_52_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1529__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_167 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_145 VGND VPWR sky130_fd_sc_hd__decap_4
X_1078_ _1078_/A _1014_/B _1078_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0995__B2 _0994_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0995__A1 _0823_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1387__A data_in[3] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1537__D _1537_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1227__A2 _1216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_370 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_42 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_53 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0986__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0986__B2 _0981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1297__A _1305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1447__D _1447_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1163__A1 _0917_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_1001_ _1537_/Q _1056_/A _1000_/Y _1001_/D _1001_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_19_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_112 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_167 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1218__A2 _1216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_318 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0977__A1 _0969_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0977__B2 _0972_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0823__B _0823_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1000__A _1539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1357__D _1356_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0716_ _0757_/B _0716_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0963__A1_N _0738_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_156 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1562__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0968__A1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0968__B2 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1393__A1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_20 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0908__B _1090_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_292 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0924__A _1155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_167 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_189 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0959__B2 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0959__A1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_300 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1081__B1 _1080_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1550_ _1550_/D _1550_/Q _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1481_ _1291_/Y _1285_/A _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_11_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0818__B _0818_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0834__A _0823_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1384__B _0935_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_clk_48_A clkbuf_4_5_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1127__A1 _1567_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0728__B _0879_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_218 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1550__D _1550_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_292 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0744__A _0743_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_67 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1063__B1 _1062_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1366__A1 _1350_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__A1 _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0919__A _1560_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_207 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0877__B1 _0892_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1460__D _1045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_0981_ _0957_/X _0981_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1054__B1 _1013_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1602_ _1235_/X _1234_/A _0928_/X _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_59_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1533_ _1533_/D _1533_/Q _0927_/X _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1464_ _1463_/Q _0806_/A _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_67_310 VGND VPWR sky130_fd_sc_hd__decap_12
X_1395_ data_in[4] _0935_/Y _1395_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0829__A _0823_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_229 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_262 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1293__B1 _1292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1379__B _0786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1045__B1 _0823_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1548__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1395__A data_in[4] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1348__A1 _1513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1545__D _1075_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__A usb_address[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_221 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0921__B _0921_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1455__D _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_1180_ _0838_/Y _1171_/X _0768_/X _1171_/X _1180_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA_clkbuf_4_11_0_clk_48_A clkbuf_3_5_0_clk_48/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1275__B1 _1269_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_284 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1562__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1027__B1 _1525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_0964_ _0740_/Y _0962_/Y _1438_/Q _0962_/Y _0964_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0895_ _1317_/A _0895_/B _0754_/D _0895_/X VGND VPWR sky130_fd_sc_hd__or3_4
X_1516_ _1516_/D _0776_/A rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_118 VGND VPWR sky130_fd_sc_hd__decap_4
X_1447_ _1447_/D _1447_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_4_81 VGND VPWR sky130_fd_sc_hd__fill_2
X_1378_ _0724_/A _1394_/D _1366_/X _1397_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_67_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_346 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0725__C _0886_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_46 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_276 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1435__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_313 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1585__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_346 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0916__B _1159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_97 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_349 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1257__B1 _1256_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_254 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1009__B1 _1008_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0932__A _0757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1024__A3 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1594__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__B1_N _1117_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1301_ _1259_/X _1300_/X _1296_/X _1301_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_1232_ _1601_/Q _1200_/A _1232_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_49_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_1163_ _0917_/X _1161_/Y _1147_/A _1162_/X _1163_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_49_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0826__B _0826_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1094_ _1090_/A _1094_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_52_327 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1003__A _1003_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1015__A3 _1014_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0947_ endpoint[0] _0945_/B _0947_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1587__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1458__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1516__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_0878_ _0855_/X _0865_/X _0870_/Y _0877_/X _0878_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__1392__B _1387_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_338 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1239__B1 _1604_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0752__A _0744_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1411__B1 _1406_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1604__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_53 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_346 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_357 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0927__A _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_327 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_371 VGND VPWR sky130_fd_sc_hd__decap_4
X_0801_ _0799_/Y _0800_/Y _0802_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1600__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1402__B1 _1381_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_261 VGND VPWR sky130_fd_sc_hd__fill_2
X_0732_ _0732_/A _0776_/B _0733_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_41_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1215_ _1212_/A _1208_/X _1214_/X _1593_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0837__A _0836_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1146_ _1145_/B usb_rst _1145_/A _1147_/C VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_37_165 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1307__A1_N _1612_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1077_ _0999_/D _1069_/X _1076_/X _1077_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_33_371 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0995__A2 _0823_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1387__B _1399_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_404 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1553__D _1553_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__A _1449_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_55 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_77 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_393 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0986__A2 _0980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1297__B _1296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1396__C1 _1395_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_264 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1163__A2 _1161_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1463__D _0798_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1000_ _1539_/Q _1000_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_19_143 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1320__C1 _0870_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_393 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0977__A2 _0971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_341 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_363 VGND VPWR sky130_fd_sc_hd__decap_3
X_0715_ _0715_/A _0715_/B _0715_/C _0757_/B VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_57_238 VGND VPWR sky130_fd_sc_hd__fill_2
X_1129_ _1102_/A _1147_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_15_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0968__A2 _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_352 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1531__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1548__D _1081_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_35 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1393__A2 _1409_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_278 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_54 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0908__C _0904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_113 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0924__B _1154_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_330 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_127 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__A2 _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_312 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_374 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1081__A1 _1078_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1458__D _1458_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0940__A setup VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1519__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1480_ _1287_/X _0708_/B _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_39_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0834__B _0834_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1011__A _1534_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0850__A _0901_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_193 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1170__A1_N _1094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1127__A2 _1123_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0744__B _0744_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_23 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1063__A1 _1539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0760__A handshake[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1366__A2 _0725_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__A2 _1114_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_39 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0919__B _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0877__B2 _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_282 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0935__A _0935_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_285 VGND VPWR sky130_fd_sc_hd__fill_2
X_0980_ _0970_/X _0980_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_120 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1054__B2 _1036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_197 VGND VPWR sky130_fd_sc_hd__decap_4
X_1601_ _1233_/X _1601_/Q _0928_/X _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1532_ _1532_/D _1532_/Q _0927_/X _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1491__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1463_ _0798_/A _1463_/Q _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_67_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_322 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0829__B _0829_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1394_ _1350_/X _0785_/X _0869_/A _1394_/D _1394_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1006__A _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0915__A1_N _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0845__A _0851_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1293__A1 _1288_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_119 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1045__B2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1045__A1 _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1395__B _0935_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1348__A2 _1346_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_322 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0739__B _0738_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1561__D _1108_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0755__A _0755_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_300 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1471__D _1191_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_325 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_399 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1275__B2 _1241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1027__B2 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1027__A1 _1020_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0963_ _0738_/Y _0962_/Y _1437_/Q _0962_/Y _1445_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0894_ _1319_/A _1340_/B _0894_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1515_ _1328_/X _1315_/A rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_4_93 VGND VPWR sky130_fd_sc_hd__decap_4
X_1446_ _0964_/X _1446_/Q _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1377_ _1400_/B _1394_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_67_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_314 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_288 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1556__D _1098_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_196 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0916__C _0916_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_87 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1257__A1 _1241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_49 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1009__A1 _1536_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1009__B2 _0841_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1466__D _1466_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_8 VGND VPWR sky130_fd_sc_hd__fill_2
X_1300_ _1300_/A _0892_/B _1299_/X _1300_/X VGND VPWR sky130_fd_sc_hd__or3_4
X_1231_ _1228_/A _1205_/X _1230_/X _1231_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_1_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_122 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_111 VGND VPWR sky130_fd_sc_hd__fill_2
X_1162_ _1159_/A _0924_/X _1162_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_358 VGND VPWR sky130_fd_sc_hd__decap_4
X_1093_ _0768_/X _1187_/C _1090_/X _0904_/A _1092_/X _1553_/D VGND VPWR sky130_fd_sc_hd__o32a_4
XFILLER_64_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1003__B _1086_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_247 VGND VPWR sky130_fd_sc_hd__decap_4
X_0946_ _0755_/A _0755_/B _0942_/X direction_in _0945_/X _0946_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_9_281 VGND VPWR sky130_fd_sc_hd__fill_2
X_0877_ _0716_/X _0872_/X _0892_/A _0876_/X _0877_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1184__B1 _1181_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1392__C _1391_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1556__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_1429_ _0986_/X data_out[2] _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_28_325 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_380 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1239__B2 _1205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1239__A1 _1214_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_391 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_372 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0752__B _0746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_23 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1411__B2 _1410_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0746__A1_N _0743_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1552__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0927__B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1104__A _1128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0989__B1 data_out[5] VGND VPWR sky130_fd_sc_hd__diode_2
X_0800_ _1466_/D _0800_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_24_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1402__A1 _1284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0731_ _0776_/A _0732_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_6_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0913__B1 _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1214_ _1593_/Q _1214_/B _1214_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1145_ _1145_/A _1145_/B usb_rst _1149_/B VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_25_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1014__A _1014_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_199 VGND VPWR sky130_fd_sc_hd__fill_2
X_1076_ _1002_/C _1064_/X _1076_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0853__A _0853_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_180 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1425__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0995__A3 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0929_ _0874_/A _1194_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1575__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1157__B1 _1155_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_114 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_34 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_158 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_11 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0_0_clk_48_A clkbuf_2_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_66 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0986__A3 _1445_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1396__B1 _1373_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0938__A _0937_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1320__B1 _1319_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1448__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_180 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0977__A3 _1524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1275__A2_N _1274_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1598__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_386 VGND VPWR sky130_fd_sc_hd__fill_2
X_0714_ _0714_/A _0715_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_217 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0848__A _0777_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_114 VGND VPWR sky130_fd_sc_hd__decap_4
X_1128_ _1128_/A _1128_/B _1128_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_65_294 VGND VPWR sky130_fd_sc_hd__fill_2
X_1059_ _1004_/X _1059_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0968__A3 _1442_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1378__B1 _1366_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1571__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1564__D _1119_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1500__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_246 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0758__A _0757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0908__D _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_77 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_131 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0924__C _1154_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_120 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_353 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0959__A3 _1435_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_324 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1081__A2 _1069_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1474__D _1271_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_253 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_191 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_286 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1202__A _1196_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1559__D _1101_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1063__A2 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_68 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0919__C _0919_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1112__A _1102_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1469__D _0766_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0951__A endpoint[2] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1493__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_1600_ _1231_/X _1600_/Q _0928_/X _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_32_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_1531_ _0995_/X _0994_/A rst_n _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1462_ rx_se0 _0798_/A _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_67_334 VGND VPWR sky130_fd_sc_hd__decap_12
X_1393_ _0785_/X _1409_/B _1386_/X _1392_/X _1422_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_67_367 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_clk_48 clkbuf_3_7_0_clk_48/X _1589_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1006__B _1006_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1293__A2 _1252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_267 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1045__A2 _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0861__A _1358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_38 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0755__B _0755_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1509__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_256 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0771__A _0771_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_109 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_323 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1107__A _1560_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_304 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_220 VGND VPWR sky130_fd_sc_hd__decap_4
X_0962_ _0961_/X _0962_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1027__A2 _1037_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_267 VGND VPWR sky130_fd_sc_hd__decap_4
X_0893_ _0775_/X _1340_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_64_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1514_ _1325_/Y _1381_/A rst_n _1514_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_4_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1017__A _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1445_ _1445_/D _1445_/Q _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_67_142 VGND VPWR sky130_fd_sc_hd__decap_4
X_1376_ _0887_/A _1400_/B _1371_/X _1374_/X _1375_/Y _1376_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_55_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0856__A _1316_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1572__D _1572_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_23 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0766__A _0766_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1257__A2 _1255_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_223 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1481__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1009__A2 _0840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_81 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1482__D _1293_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_7 VGND VPWR sky130_fd_sc_hd__decap_4
X_1230_ _1600_/Q _1222_/B _1230_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_1_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_101 VGND VPWR sky130_fd_sc_hd__fill_1
X_1161_ _1160_/X _1161_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_64_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VPWR sky130_fd_sc_hd__fill_2
X_1092_ _1095_/A _1092_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1003__C _1550_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_215 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1300__A _1300_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0945_ _0754_/B _0945_/B _0945_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_293 VGND VPWR sky130_fd_sc_hd__fill_2
X_0876_ _1187_/A tx_en _0876_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1184__A1 _1095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_48_A clkbuf_3_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1428_ _0985_/X data_out[1] _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1061__A1_N _1016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_1359_ _0886_/A _1354_/X _1355_/X _1357_/X _1358_/X _1359_/X VGND VPWR sky130_fd_sc_hd__a2111o_4
XANTENNA__1525__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_359 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1239__A2 _1238_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_36 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_204 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0752__C _0749_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1567__D _1128_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_167 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1104__B _1104_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0989__B2 _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0989__A1 _0901_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_351 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1120__A _0920_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_384 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1477__D _1279_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0730_ _1317_/A _0895_/B _0754_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1402__A2 _1409_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0913__A1 _1102_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1213_ _1591_/Q _1208_/X _1212_/X _1213_/X VGND VPWR sky130_fd_sc_hd__a21o_4
Xclkbuf_4_2_0_clk_48 clkbuf_4_3_0_clk_48/A _1443_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_27_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_123 VGND VPWR sky130_fd_sc_hd__fill_2
X_1144_ _1158_/A _1144_/B _1143_/Y _1144_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_1_62 VGND VPWR sky130_fd_sc_hd__decap_4
X_1075_ _1072_/A _1069_/X _1074_/X _1075_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1014__B _1014_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_362 VGND VPWR sky130_fd_sc_hd__decap_4
X_0928_ rst_n tx_en _0928_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0859_ _0858_/X _1413_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1157__A1 _1155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1205__A _1205_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_318 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1093__B1 _0904_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0840__B1 _1461_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1396__A1 _1423_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1320__A1 _1315_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_126 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0831__B1 _0829_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_398 VGND VPWR sky130_fd_sc_hd__fill_2
X_0713_ _0713_/A _1300_/A _0714_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_1127_ _1567_/Q _1123_/X _1130_/B _1128_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XANTENNA__1311__A1 _1309_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0864__A _0861_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_148 VGND VPWR sky130_fd_sc_hd__fill_2
X_1058_ _1056_/Y _1036_/X _1537_/Q _1057_/X _1538_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1075__B1 _1074_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_310 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1542__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1378__A1 _0724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_12 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1580__D _1173_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_240 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0774__A _1513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_159 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_132 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1066__B1 _1065_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_118 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_192 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0949__A endpoint[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_218 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1490__D _0878_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1565__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_265 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1537__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0804__B1 _0803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_48_A clk_48 VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_94 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0859__A _0858_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_254 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1202__B _1202_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1575__D _1575_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1438__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0769__A _1495_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0919__D _0919_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_99 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1588__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1287__B1 _0708_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_232 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0951__B _0945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_173 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1485__D _0847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1211__B1 _1591_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_1530_ _1530_/D _0791_/A rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1461_ _1180_/X _1461_/Q _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1392_ _0886_/A _1387_/X _1391_/X _1392_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_67_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1278__B1 _0707_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1303__A _1303_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0755__C _1329_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_46 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0771__B _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1107__B _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_349 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1123__A _0921_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_clk_48_A clkbuf_4_5_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0962__A _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_246 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1027__A3 _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0961_ _0957_/X _0961_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0847__B1_N _0846_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1603__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0892_ _0892_/A _0892_/B _0892_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_57_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1513_ _1513_/D _1513_/Q rst_n _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1444_ _0960_/X _1444_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1375_ _1409_/A _1372_/X _0935_/Y _1375_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0856__B _0856_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_371 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_213 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0872__A _0769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_257 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1208__A _1205_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_132 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0766__B _0766_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_305 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1244__A1_N _1250_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0957__A _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_110 VGND VPWR sky130_fd_sc_hd__fill_2
X_1160_ _1160_/A _1160_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_37_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_1091_ _1090_/A _1095_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_64_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_371 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1003__D _1003_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_363 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1300__B _0892_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0944_ _0755_/A _0941_/X _0943_/X _0944_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1405__B1 _1284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0875_ _0874_/X tx_en VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1184__A2 _1183_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1427_ _1427_/D data_out[0] _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0867__A _0760_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_1358_ _1358_/A _0775_/X _1358_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1289_ _1406_/A _1289_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1058__A2_N _1036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1565__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0752__D _0751_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_69 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_10_0_clk_48_A clkbuf_3_5_0_clk_48/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1583__D _1177_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0777__A _0777_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1332__C1 _1331_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0989__A2 _0970_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1401__A _0887_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1120__B _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_70 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_81 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1493__D _1493_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0913__A2 _0824_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1212_ _1212_/A _1214_/B _1212_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_65_400 VGND VPWR sky130_fd_sc_hd__decap_6
X_1143_ _1143_/A _1139_/X _1143_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_1_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_157 VGND VPWR sky130_fd_sc_hd__fill_2
X_1074_ _0999_/D _1064_/X _1074_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1014__C _1013_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_168 VGND VPWR sky130_fd_sc_hd__fill_2
X_0927_ _0885_/A rst_n _0927_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0858_ _1528_/Q _0994_/B _0858_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1157__A2 _1156_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0789_ _0788_/X _0789_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1471__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_48 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_127 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1578__D _1578_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_374 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1093__A1 _0768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1093__B2 _1092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0840__A1 _0838_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0840__B2 _1187_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1396__A2 _1394_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_70 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1487__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1320__A2 _0794_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1131__A _1131_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_322 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1488__D _1488_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0970__A _1413_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0831__B2 _0830_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0712_ _0712_/A _0712_/B _1612_/Q _1300_/A VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__1494__CLK _1514_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1306__A _1304_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_252 VGND VPWR sky130_fd_sc_hd__fill_2
X_1126_ _0922_/D _0925_/Y _1130_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_53_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1311__A2 _1300_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0864__B _0864_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1057_ _0994_/B _1057_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1075__A1 _1072_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_119 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0880__A _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1378__A2 _1394_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1216__A _1205_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_24 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1580__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0774__B _0773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_300 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1066__A1 _1540_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_322 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_304 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_71 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0949__B _0945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1126__A _0922_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_252 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0804__A1 _0797_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1036__A _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0875__A _0874_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1109_ _0919_/C _1109_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_53_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1591__D _1591_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1543__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0785__A _1357_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1287__B2 _1240_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_145 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1211__A1 _1214_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1211__B2 _1205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_1460_ _1045_/X _0823_/A _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1391_ _0758_/Y _1391_/B _1391_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1532__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_358 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1278__A1 _1388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1303__B _1298_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1519__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_314 VGND VPWR sky130_fd_sc_hd__fill_2
X_1589_ _1589_/D _1589_/Q _0928_/X _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_58_369 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_236 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0771__C _1509_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1586__D _1182_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1555__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0952__B1 _0951_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1107__C _1150_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_358 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1123__B _1150_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_288 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_299 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1115__B1_N _1114_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0960_ _0855_/X _0955_/X _1436_/Q _1444_/Q _0958_/X _0960_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_32_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1496__D _1360_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0891_ _0890_/Y _0891_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1512_ _1512_/D _1512_/Q rst_n _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1612__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_1443_ _0959_/X _1443_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0943__B1 _0940_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_85 VGND VPWR sky130_fd_sc_hd__decap_3
X_1374_ _1420_/Q _1373_/Y _1374_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_328 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1428__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_236 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0872__B _1409_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1578__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1224__A _1597_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_24 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1178__B1 _1583_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_184 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0957__B _0957_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1134__A _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_199 VGND VPWR sky130_fd_sc_hd__decap_3
X_1090_ _1090_/A _1090_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_64_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_331 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1300__C _1299_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0943_ _0895_/B _0942_/X _0940_/Y _0943_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1405__B2 _1410_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_0874_ _0874_/A _0874_/B _0874_/C _0874_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1169__B1 _1158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1309__A _1309_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1426_ _1412_/X _1406_/A _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0867__B _0867_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1007__B1_N _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1357_ _1350_/X _1357_/B _1329_/A _1356_/X _1357_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_55_147 VGND VPWR sky130_fd_sc_hd__fill_2
X_1288_ _1482_/Q _1288_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0883__A tx_en VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_16 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_228 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1219__A _1200_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__B _0777_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1332__B1 _1330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0793__A _0732_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_180 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0989__A3 _0744_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1401__B _1399_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1120__C _0920_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1103__A2_N usb_rst VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1129__A _1102_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1211_ _1214_/B _1210_/X _1591_/Q _1205_/X _1591_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_37_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1323__B1 _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1142_ _1143_/A _1139_/X _1144_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_1_53 VGND VPWR sky130_fd_sc_hd__fill_2
X_1073_ _0999_/B _1069_/X _1072_/X _1073_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1014__D _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_353 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_397 VGND VPWR sky130_fd_sc_hd__fill_2
X_0926_ _0925_/Y usb_rst VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1039__A _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0857_ _0816_/X _0994_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_0788_ _1324_/A _1315_/A _0788_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_1409_ _1409_/A _1409_/B _1408_/X _1409_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_68_261 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1314__B1 _0935_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1093__A2 _1187_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0840__A2 _0768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1594__D _1218_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_268 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0788__A _1324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_250 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_353 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_397 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_334 VGND VPWR sky130_fd_sc_hd__fill_2
X_0711_ _1305_/A _0712_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1306__B _1306_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_242 VGND VPWR sky130_fd_sc_hd__fill_2
X_1125_ _1128_/A _1125_/B _1125_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__1322__A _0869_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_18 VGND VPWR sky130_fd_sc_hd__fill_2
X_1056_ _1056_/A _1056_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_18_180 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1075__A2 _1069_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0880__B _0783_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_367 VGND VPWR sky130_fd_sc_hd__decap_4
X_0909_ _0768_/X _1187_/C _0909_/C _0908_/X _0909_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_0_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_36 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_253 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1232__A _1601_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1589__D _1589_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1066__A2 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_172 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_334 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_378 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_316 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1126__B _0925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_404 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_275 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1142__A _1143_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1499__D _0952_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0981__A _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0804__A2 _0802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1461__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1317__A _1317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_286 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_1108_ _1105_/X _1107_/Y _1187_/C _1108_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_53_278 VGND VPWR sky130_fd_sc_hd__fill_2
X_1039_ _0994_/B _1039_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0891__A _0890_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_297 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1484__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_267 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_289 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1089__A1_N _1016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1211__A2 _1210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1137__A _1137_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_1390_ _1388_/Y _1362_/X _1389_/X _1391_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_67_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1278__A2 _1273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1303__C _1302_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_278 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_1588_ _0768_/X _1588_/Q rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__0886__A _0886_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1559__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_267 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0952__A1 _1436_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_0890_ _0777_/A _0890_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_43_92 VGND VPWR sky130_fd_sc_hd__fill_2
X_1511_ _1345_/X _0772_/C rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1442_ _0983_/X _1442_/Q _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0943__A1 _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_123 VGND VPWR sky130_fd_sc_hd__fill_2
X_1373_ _0725_/B _1372_/X _1373_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_67_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1330__A _1330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0790__A1_N _0887_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_119 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1224__B _1222_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_329 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_215 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1240__A _0715_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1597__D _1225_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1522__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1178__B2 _1171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1415__A _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_123 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1134__B _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_126 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1150__A _1154_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_0942_ _0938_/X _0942_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_285 VGND VPWR sky130_fd_sc_hd__fill_2
X_0873_ _0873_/A _0874_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_62_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1169__A1 _0916_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1425_ _1425_/D _1425_/Q _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1356_ _0777_/A _0862_/A _1492_/Q _1356_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_28_329 VGND VPWR sky130_fd_sc_hd__fill_2
X_1287_ _1272_/X _1286_/X _0708_/B _1240_/X _1287_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_362 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_395 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1545__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_343 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_49 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1574__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1411__A1_N _0769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_58 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1503__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1332__A1 _0771_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0793__B _1316_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1096__B1 _1554_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_192 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1401__C _1401_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1120__D _0925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_71 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1145__A _1145_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1210_ _1207_/A _1204_/Y _1207_/Y _1204_/A _1210_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_1141_ _0918_/A _1143_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1323__B2 _1322_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1323__A1 _0861_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1568__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1072_ _1072_/A _1064_/X _1072_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1087__B1 _1550_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1287__A2_N _1286_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_184 VGND VPWR sky130_fd_sc_hd__decap_4
X_0925_ _0917_/X _0924_/X _0925_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0856_ _1316_/B _0856_/B _0856_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0787_ _1381_/A _1324_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_1408_ _1289_/Y _1381_/X _1408_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_56_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1314__A1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_284 VGND VPWR sky130_fd_sc_hd__fill_2
X_1339_ _0772_/A _0772_/B _1339_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0894__A _1319_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_38 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_343 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_365 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1093__A3 _1090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_37 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_195 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_203 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_41 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0788__B _1315_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1589__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_1_0_clk_48_A clkbuf_3_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_376 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_195 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_368 VGND VPWR sky130_fd_sc_hd__fill_2
X_0710_ _0709_/X _0713_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_51_70 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1496__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0979__A _1187_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1306__C _1301_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_210 VGND VPWR sky130_fd_sc_hd__fill_2
X_1124_ _1566_/Q _1120_/X _1123_/X _1125_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_65_298 VGND VPWR sky130_fd_sc_hd__decap_3
X_1055_ _1046_/X _1004_/X _1537_/Q _1016_/X _1537_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1322__B _1358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0807__B1 _0806_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_29 VGND VPWR sky130_fd_sc_hd__decap_4
X_0908_ _1557_/Q _1090_/A _0904_/X _0907_/X _0908_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0889__A _0789_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0839_ _0768_/X _1187_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_0_206 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1299__B1 _1604_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1232__B _1200_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_151 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_328 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_2_0_clk_48 clkbuf_3_3_0_clk_48/A clkbuf_4_5_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1223__B1 _1222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_40 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0799__A _1466_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_202 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1142__B _1139_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_81 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1606__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_184 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1606__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_350 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1317__B _0755_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1333__A _0771_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_1107_ _1560_/Q _0919_/B _1150_/B _1107_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_53_268 VGND VPWR sky130_fd_sc_hd__fill_2
X_1038_ _1036_/X _0827_/B _1037_/X _1038_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_21_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1243__A _0874_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1418__A _1605_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1137__B _1137_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0992__A _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_227 VGND VPWR sky130_fd_sc_hd__fill_2
X_1587_ _1184_/X _1587_/Q rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_37_28 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1528__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_249 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0952__A2 _0942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1451__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_327 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0911__A1_N _0818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1417__B1 _1296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1148__A _1573_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1510_ _1510_/D _0772_/A rst_n _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_4_150 VGND VPWR sky130_fd_sc_hd__decap_3
X_1441_ _0982_/X _1441_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_4_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0943__A2 _0942_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1372_ _1409_/A _0889_/Y _0769_/Y _1372_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_67_146 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_5_0_clk_48 clkbuf_4_5_0_clk_48/A _1567_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_293 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1474__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_113 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_341 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_374 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_227 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_153 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1415__B _1415_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_146 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_105 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1134__C _0922_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_71 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1150__B _1150_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_208 VGND VPWR sky130_fd_sc_hd__fill_2
X_0941_ _0895_/B _0945_/B _0940_/Y _0941_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_9_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_293 VGND VPWR sky130_fd_sc_hd__fill_2
X_0872_ _0769_/Y _1409_/A _0872_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1497__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1169__A2 _1165_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1424_ _1424_/D _1424_/Q _1514_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1355_ _1319_/A _1318_/A _1355_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_138 VGND VPWR sky130_fd_sc_hd__fill_2
X_1286_ _1284_/Y _1247_/D _1285_/Y _1286_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1341__A _1340_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_193 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_333 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_3_0_clk_48_A clkbuf_4_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1332__A2 _1340_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_300 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1096__B2 _1095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1096__A1 _0904_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_322 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_234 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1549__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_8 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1145__B _1145_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_81 VGND VPWR sky130_fd_sc_hd__fill_2
X_1140_ _1137_/X _1139_/X _1158_/A _1570_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1323__A2 _0778_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1161__A _1160_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1071_ _0999_/C _1069_/X _1070_/X _1071_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_1_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_341 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1087__B2 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_141 VGND VPWR sky130_fd_sc_hd__fill_2
X_0924_ _1155_/A _1154_/A _1154_/B _0924_/X VGND VPWR sky130_fd_sc_hd__or3_4
X_0855_ _1187_/A _0855_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0786_ _0722_/X _0786_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1336__A _0771_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_230 VGND VPWR sky130_fd_sc_hd__decap_12
X_1407_ _1389_/X _1406_/X _1399_/B data_in[7] _0758_/Y _1407_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1512__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1314__A2 _1313_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1338_ _0775_/X _1337_/Y _1330_/X _1509_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_28_127 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0894__B _1340_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1269_ _1269_/A _1269_/B _1269_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_28 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_333 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1246__A _0715_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_108 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_141 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_174 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1156__A _0917_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1535__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_266 VGND VPWR sky130_fd_sc_hd__fill_2
X_1123_ _0921_/B _1150_/B _1123_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_1054_ _1008_/Y _1036_/X _1013_/C _1036_/X _1054_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__0807__A1 _0797_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_152 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_336 VGND VPWR sky130_fd_sc_hd__decap_3
X_0907_ _1555_/Q _0905_/Y _0906_/Y _0907_/D _0907_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1532__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1595__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0991__B1 data_out[7] VGND VPWR sky130_fd_sc_hd__diode_2
X_0838_ _1461_/Q _0838_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0769_ _1495_/Q _0769_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_0_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_16 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1299__B2 _1196_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_406 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_303 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_196 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1223__A1 _1595_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_391 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1558__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0982__B1 _1441_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_52 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0734__B1 usb_address[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_269 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0973__B1 _1435_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1317__C _0890_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_211 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1333__B _1340_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1106_ _0925_/Y _1150_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_53_214 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_1037_ _1037_/A _0912_/X _1037_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_42_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0964__B1 _1438_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1243__B _0715_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1178__A2_N _1171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0946__B1 direction_in VGND VPWR sky130_fd_sc_hd__diode_2
X_1586_ _1182_/Y _1183_/B rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_328 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1344__A _0772_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1568__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1254__A _0874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_309 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1417__A1 _1606_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_50 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1209__A1_N _1207_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1440_ _0978_/X _1440_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_4_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_195 VGND VPWR sky130_fd_sc_hd__fill_2
X_1371_ data_in[1] _1399_/B _1371_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1164__A _0916_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_99 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1353__B1 _0764_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_91 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1105__B1 _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_375 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1339__A _0772_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__A2_N _1004_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1569_ _1135_/X _0922_/B rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1074__A _0999_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_353 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_206 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1249__A _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1180__A1_N _0838_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1415__C _1415_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1134__D _1150_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_389 VGND VPWR sky130_fd_sc_hd__fill_2
X_0940_ setup _0940_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1159__A _1159_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0871_ _1357_/B _1409_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0998__A _0997_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1423_ _1396_/X _1423_/Q _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_48_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1326__B1 _1327_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1354_ data_in_valid _0887_/D _0757_/B _1354_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_55_106 VGND VPWR sky130_fd_sc_hd__decap_4
X_1285_ _1285_/A _1285_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_48_180 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_161 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_367 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1441__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1069__A _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1591__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_128 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_353 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1583__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1096__A2 _1094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1512__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_74 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_40 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1145__C usb_rst VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_23 VGND VPWR sky130_fd_sc_hd__fill_2
X_1070_ _0999_/B _1064_/X _1070_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_65_81 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_70 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_120 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_323 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1464__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_0923_ _1573_/Q _1145_/A _1145_/B _1154_/B VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1087__A1_N _1086_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0854_ _0885_/A _0818_/X _0853_/Y _1487_/D VGND VPWR sky130_fd_sc_hd__a21o_4
X_0785_ _1357_/B _0785_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1336__B _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1406_ _1406_/A _1362_/X _1406_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_253 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_242 VGND VPWR sky130_fd_sc_hd__decap_6
X_1337_ _1335_/Y _1336_/Y _0772_/B _1337_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_68_275 VGND VPWR sky130_fd_sc_hd__decap_4
X_1268_ _1247_/D _1269_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1502__D _0944_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1199_ _1205_/A _1200_/A VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_142 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1262__A _1250_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1487__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_326 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1172__A _0813_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_245 VGND VPWR sky130_fd_sc_hd__decap_4
X_1122_ _1128_/A _1122_/B _1122_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_65_278 VGND VPWR sky130_fd_sc_hd__decap_3
X_1053_ _1014_/A _1046_/X _1013_/C _1046_/X _1053_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0807__A2 _0803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_304 VGND VPWR sky130_fd_sc_hd__fill_1
X_0906_ _0906_/A _0906_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0991__A1 _0901_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0837_ _0836_/X _0837_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0768_ _0767_/X _0768_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0991__B2 _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1082__A _1002_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_223 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_109 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_115 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_326 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_308 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1223__A2 _1216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0982__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0982__B2 _0981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0734__B2 _1443_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_267 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0741__A1_N usb_address[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_164 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1502__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_189 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1167__A _0916_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0973__A1 _0969_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0973__B2 _0972_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_99 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1317__D _1317_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1333__C _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_234 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_1105_ _1560_/Q usb_rst _0919_/B _1105_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_38_267 VGND VPWR sky130_fd_sc_hd__fill_2
X_1036_ _0992_/X _1036_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_61_292 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0964__B2 _0962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1525__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1127__B1_N _1130_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1600__D _1231_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0946__B2 _0945_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0946__A1 _0755_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1585_ _1179_/X _0814_/C rst_n _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_318 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1344__B _1342_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_215 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1548__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0882__B1 _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1510__D _1510_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1019_ _1528_/Q _1016_/X _1018_/X _1019_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_34_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_281 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1254__B _1252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_373 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1270__A _1363_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1420__D _1376_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1417__A2 _1605_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1050__B1 _1533_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_23 VGND VPWR sky130_fd_sc_hd__fill_2
X_1370_ _1369_/X _1400_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_70 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1164__B _1160_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1353__A1 _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1105__A1 _1560_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1339__B _0772_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1041__B1 _0836_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1355__A _1319_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1568_ _1568_/D _0922_/A rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1074__B _1064_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1499_ _0952_/X endpoint[2] rst_n _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1505__D _1353_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_321 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1090__A _1090_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1280__B1 _0707_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1249__B _0715_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1032__B1 _1317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1265__A _0715_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1099__B1 _1557_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_273 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1271__B1 _1201_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1159__B _0924_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_277 VGND VPWR sky130_fd_sc_hd__fill_2
X_0870_ data_in_valid _0887_/D _0870_/C _0870_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__1023__B1 _1521_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1422_ _1422_/D _1388_/A _1514_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1175__A _0813_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1326__A1 _0869_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1353_ _0716_/X _1352_/X _0764_/X _1353_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_1284_ _1425_/Q _1284_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_36_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_398 VGND VPWR sky130_fd_sc_hd__fill_2
X_0999_ _1540_/Q _0999_/B _0999_/C _0999_/D _1005_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_39_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_184 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1253__B1 _1252_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_254 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_151 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1609__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_154 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1054__A2_N _1036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_379 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1244__B1 _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0922_ _0922_/A _0922_/B _0922_/C _0922_/D _1145_/B VGND VPWR sky130_fd_sc_hd__or4_4
X_0853_ _0853_/A _0853_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0802__A _0798_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_0784_ _0769_/Y _0887_/B _0783_/X _1495_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1405_ _1401_/X _1404_/X _1284_/Y _1410_/B _1425_/D VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
X_1336_ _0771_/A _0771_/B _1336_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_1267_ _1272_/A _1267_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_1198_ _1473_/Q _1196_/Y _1252_/B _1205_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_18 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1235__B1 _1234_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__A _0712_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0831__A2_N _0830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_298 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1262__B _1245_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_357 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_305 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1172__B _1090_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_235 VGND VPWR sky130_fd_sc_hd__decap_4
X_1121_ _0920_/A _1117_/X _1120_/X _1122_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XANTENNA__1431__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1603__D _1237_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_1052_ _1046_/X _1050_/X _1051_/X _1052_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_18_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1581__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_176 VGND VPWR sky130_fd_sc_hd__decap_3
X_0905_ _1556_/Q _0905_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0991__A2 _0970_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0836_ _0821_/Y _0836_/B _0836_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0767_ _0766_/A _0766_/B _1467_/Q _0766_/X _0767_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1363__A _1363_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1153__C1 _1152_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1082__B _1014_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1513__D _1513_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1319_ _1319_/A _1318_/Y _1319_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_56_257 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0707__A _0707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_143 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_176 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_349 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0982__A2 _0980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_98 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1454__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1273__A _1269_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1423__D _1396_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_73 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_168 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_371 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_56 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1167__B _1160_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0973__A2 _0971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1183__A _1587_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__C1 _1137_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1104_ _1128_/A _1104_/B _1104_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_1035_ _0826_/B _0992_/X _1034_/X _0840_/X _1035_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_21_102 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1358__A _1358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1508__D _1334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1477__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0819_ _0901_/B _0846_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_3_0_0_clk_48_A clkbuf_3_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_268 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_87 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1268__A _1247_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_97 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_293 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0946__A2 _0755_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__A _1587_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1584_ _1178_/X _0811_/A rst_n _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xclkbuf_2_2_0_clk_48 clkbuf_2_3_0_clk_48/A clkbuf_3_5_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_26_238 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0882__A1 _0879_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1018_ _1018_/A _1018_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xclkbuf_4_10_0_clk_48 clkbuf_3_5_0_clk_48/X _1611_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0720__A _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1577__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1506__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1254__C _0874_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_216 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1270__B _1247_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_293 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1050__A1 _1048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1050__B2 _1010_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1353__A2 _1352_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1105__A2 usb_rst VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_385 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1611__D _1306_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_260 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_219 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_399 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0805__A _1466_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1041__A1 _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1041__B2 _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1567_ _1128_/Y _1567_/Q rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1355__B _1318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1515__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1498_ _1498_/D endpoint[1] rst_n _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1371__A data_in[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1521__D _1521_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_219 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1538__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0715__A _0715_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1280__A1 _1423_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1032__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1032__B2 _0853_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1265__B _0892_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_74 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1099__B2 _1095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1099__A1 _1556_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1431__D _1431_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_252 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1271__A1 _1267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1271__B2 _1240_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_245 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1023__A1 _1020_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1499__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1023__B2 _1021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1538__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1421_ _1385_/X _1421_/Q _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1175__B _1090_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__B1 _0755_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1606__D _1417_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1326__A2 _0725_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1352_ _1350_/X _1351_/X _0759_/X _1185_/B _1352_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_1283_ _1272_/X _1282_/Y _0707_/C _1240_/X _1283_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_152 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1299__A2_N _1196_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_358 VGND VPWR sky130_fd_sc_hd__fill_2
X_0998_ _0997_/X _0998_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1237__A2_N _1208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1516__D _1516_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_108 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0828__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_196 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_347 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1253__A1 _1241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_215 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_clk_48 clkbuf_3_5_0_clk_48/A clkbuf_3_5_0_clk_48/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_288 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1521__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0764__B1 _0886_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1426__D _1412_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_69 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_344 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_358 VGND VPWR sky130_fd_sc_hd__fill_2
X_0921_ _1567_/Q _0921_/B _0922_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_60_199 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1244__B2 _1250_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_391 VGND VPWR sky130_fd_sc_hd__fill_2
X_0852_ _0851_/X _0853_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1609__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0802__B _0802_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0783_ _1327_/B _0783_/B _0783_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1186__A _1186_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_200 VGND VPWR sky130_fd_sc_hd__fill_2
X_1404_ _0785_/X _1402_/Y _1410_/B _1403_/X _1404_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_1335_ _1509_/Q _1335_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_56_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1180__B1 _0768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_299 VGND VPWR sky130_fd_sc_hd__fill_2
X_1266_ _1265_/X _1272_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_141 VGND VPWR sky130_fd_sc_hd__fill_2
X_1197_ _0715_/C _1252_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1235__A1 _1601_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_391 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0712__B _0712_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_45 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0746__B1 _0745_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_336 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0903__A _1554_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0985__B1 data_out[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_214 VGND VPWR sky130_fd_sc_hd__fill_2
X_1120_ _0920_/A _0920_/B _0920_/C _0925_/Y _1120_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_38_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_1051_ _1014_/A _0992_/X _1051_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_4_2_0_clk_48_A clkbuf_4_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_391 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0813__A _0813_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0904_ _0904_/A _0904_/B _0904_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0976__B1 _1438_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0835_ _0835_/A _0835_/B _0843_/C VGND VPWR sky130_fd_sc_hd__xnor2_4
X_0766_ _0766_/A _0766_/B _0766_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0991__A3 _1450_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1363__B _1362_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1153__B1 _1147_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0900__B1 _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1318_ _1318_/A _1318_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_2_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_1249_ _0759_/X _0715_/B _1254_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_64_280 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0707__B _0707_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_199 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0723__A _0722_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__B1 _1441_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_33 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0982__A3 _1526_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1053__A2_N _1046_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__B1_N _0748_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_214 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_291 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0973__A3 _1520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1383__B1 _1382_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1183__B _1183_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__B1 _1147_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0808__A _0808_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1103_ _1560_/Q usb_rst _1560_/Q usb_rst _1104_/B VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
Xclkbuf_4_8_0_clk_48 clkbuf_4_9_0_clk_48/A _1421_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1034_ _1014_/B _1034_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_61_261 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_136 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1358__B _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0818_ _1102_/A _0818_/B _0818_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_0749_ usb_address[6] _0747_/Y _0748_/X _0749_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__1374__A _1420_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1524__D _1026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_236 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0718__A _0717_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_22 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_65 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1421__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1284__A _1425_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1488__SET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1571__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1434__D _1434_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_209 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1609__D _1609_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_162 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0946__A3 _0942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1356__B1 _1492_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1194__A _1250_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1583_ _1177_/X _1583_/Q rst_n _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__0810__B _1183_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1108__B1 _1187_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0882__A2 _0881_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1017_ _0998_/X _1018_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1444__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1369__A _0758_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1519__D _1519_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1594__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1347__B1 _1512_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1254__D _1254_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_272 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_220 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_75 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1429__D _0986_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1050__A2 _1009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1338__B1 _1330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_69 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_320 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1467__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_209 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0877__A1_N _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__B _1466_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1189__A _0718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_264 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1041__A2 _0835_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__A _0994_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1566_ _1125_/Y _1566_/Q rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_128 VGND VPWR sky130_fd_sc_hd__fill_2
X_1497_ _1497_/D endpoint[0] rst_n _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1371__B _1399_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_389 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0715__B _0715_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1280__A2 _1273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1032__A2 _0853_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1405__A2_N _1404_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1099__A2 _1094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_74 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0906__A _0906_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_359 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1271__A2 _1269_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_235 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1023__A2 _0829_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__A1 _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1420_ _1376_/X _1420_/Q _1514_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0782__B2 _1389_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_404 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1544__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1351_ _0759_/X _0789_/X _0785_/X _1351_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_1282_ _1424_/Q _1273_/X _0708_/B _1282_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_63_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_356 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_197 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_175 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0816__A _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0997_ _0891_/X _0816_/X _0846_/C _0997_/X VGND VPWR sky130_fd_sc_hd__or3_4
X_1549_ _1549_/D _1002_/D _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1382__A _1357_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1532__D _1532_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_131 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0828__A2 _0827_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_367 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0726__A _1317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1253__A2 _1251_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_370 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0764__A1 _0758_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1561__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1442__D _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_348 VGND VPWR sky130_fd_sc_hd__decap_3
X_0920_ _0920_/A _0920_/B _0920_/C _1566_/Q _0921_/B VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1505__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0851_ _0846_/A _0816_/X _0846_/C _0851_/D _0851_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0782_ _0895_/B data_toggle _0755_/B _1389_/D _0783_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_5_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_212 VGND VPWR sky130_fd_sc_hd__decap_4
X_1403_ _1425_/Q _0786_/Y _1350_/X _1403_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_1334_ _0771_/A _0771_/B _1330_/X _1333_/Y _1334_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_1265_ _0715_/C _0892_/B _1265_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1180__B2 _1171_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1196_ _1196_/A _1196_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_24_304 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_167 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1235__A2 _1205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_370 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1377__A _1400_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__C _1612_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0746__B2 _1444_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1527__D _1527_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_234 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1590__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1528__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_329 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0985__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1283__A2_N _1282_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0985__B2 _0981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1437__D _0975_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_226 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_131 VGND VPWR sky130_fd_sc_hd__fill_2
X_1050_ _1048_/Y _1009_/X _1533_/Q _1010_/Y _1050_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_33_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0813__B _0813_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0903_ _1554_/Q _0904_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0976__A1 _0969_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0976__B2 _0972_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0834_ _0823_/B _0834_/B _0835_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1197__A _0715_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0765_ _0725_/X _0755_/X _0764_/X _0765_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1363__C _0758_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1153__A1 _1154_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1600__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0900__B2 _0899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0900__A1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1317_ _1317_/A _0755_/B _0890_/Y _1317_/D _1318_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_1248_ _1250_/A _1245_/X _0874_/C _1248_/X VGND VPWR sky130_fd_sc_hd__and3_4
XPHY_107 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0707__C _0707_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_123 VGND VPWR sky130_fd_sc_hd__fill_2
X_1179_ _0811_/A _1090_/X _0814_/C _1092_/X _1179_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_129 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_318 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0967__B2 _0962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_384 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_56 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_207 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_86 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0914__A _0910_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1383__A1 _1421_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__A1 _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_1102_ _1102_/A _1128_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0808__B _0808_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1033_ _0837_/X _0853_/A _0755_/B _0853_/Y _1519_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_61_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0824__A _1187_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__B1 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0817_ _0816_/X _0818_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1359__D1 _1358_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0748_ usb_address[6] _0747_/Y _0748_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1374__B _1373_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1540__D _1540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_11 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0967__A2_N _0962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0909__A _0768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_96 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_218 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1450__D _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_273 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1053__B1 _1013_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_196 VGND VPWR sky130_fd_sc_hd__decap_4
X_1582_ _1582_/D _0813_/C rst_n _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1356__A1 _0777_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1194__B _1194_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1108__A1 _1105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0819__A _0901_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_229 VGND VPWR sky130_fd_sc_hd__decap_3
X_1016_ _0912_/X _1016_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1292__B1 _0715_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1369__B _1362_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1044__B1 _0832_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1347__A1 _0772_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1535__D _1053_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0729__A _0755_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_207 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1586__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1283__B1 _0707_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1515__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1035__B1 _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1295__A _0713_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1338__A1 _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_166 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1445__D _1445_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1274__B1 _0707_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_284 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0805__C _0798_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1026__B1 _1524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1122_/Y _0920_/A rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1496_ _1360_/X transaction_active rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_39_321 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_379 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1561__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0715__C _0715_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_327 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_305 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1256__B1 _1250_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1271__A3 _1270_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0922__A _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_9 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1023__A3 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__A2 data_toggle VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1350_ _1495_/Q _1350_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1434__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1281_ _1272_/X _1280_/Y _0707_/D _1240_/X _1281_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_313 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1584__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0832__A _0821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0996_ _0901_/B _0851_/D _0846_/C _0993_/X _0996_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_8_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_405 VGND VPWR sky130_fd_sc_hd__fill_2
X_1548_ _1081_/X _1003_/A _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1382__B _1381_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1479_ _1283_/X _0707_/C _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_27_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1238__B1 _1236_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0742__A _0736_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1550__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1457__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0764__A2 _0763_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0917__A _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_49 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1530__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1229__B1 _1228_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_390 VGND VPWR sky130_fd_sc_hd__fill_2
X_0850_ _0901_/A _0885_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0781_ data_toggle _1389_/D VGND VPWR sky130_fd_sc_hd__inv_8
X_1402_ _1284_/Y _1409_/B _1381_/X _1402_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_39_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1333_ _0771_/A _1340_/B _0771_/B _1333_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_1264_ _1241_/X _1261_/X _1263_/X _1609_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0827__A _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1195_ _1194_/X _1196_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_165 VGND VPWR sky130_fd_sc_hd__fill_2
X_0979_ _1187_/A _0979_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_224 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1543__D _1071_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_34 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0737__A _0856_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_371 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0985__A2 _0980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_264 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1453__D _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0813__C _0813_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0902_ _0810_/X _1090_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0976__A2 _0971_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0833_ _0833_/A _0835_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0764_ _0758_/Y _0763_/X _0886_/A _0764_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1153__A2 _1154_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1316_ _0776_/A _1316_/B _1317_/D VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0900__A2 _0889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_249 VGND VPWR sky130_fd_sc_hd__fill_2
X_1247_ _0874_/C _0874_/A _1245_/X _1247_/D _1247_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_1178_ _0811_/Y _1171_/X _1583_/Q _1171_/X _1178_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0707__D _0707_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_113 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_119 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_168 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1388__A _1388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_330 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1538__D _1538_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1298__A _0712_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1448__D _0966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0930__A _1194_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1383__A2 _1409_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1124__B1_N _1123_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1135__A2 _1131_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_249 VGND VPWR sky130_fd_sc_hd__fill_2
X_1101_ _0906_/A _1090_/X _0907_/D _1092_/X _1101_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_53_219 VGND VPWR sky130_fd_sc_hd__decap_4
X_1032_ _0827_/A _0853_/A _1317_/A _0853_/Y _1518_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0824__B _0824_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1001__A _1537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__A1 _0999_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0816_ _0815_/X _0816_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1359__C1 _1357_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0747_ _1449_/Q _0747_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1518__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0750__A usb_address[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_20 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0909__B _1187_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0925__A _0917_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_403 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1053__B2 _1046_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_175 VGND VPWR sky130_fd_sc_hd__fill_2
X_1581_ _1174_/X _1581_/Q rst_n _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1356__A2 _0862_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1108__A2 _1107_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_322 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_366 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_355 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_282 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0835__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1015_ _1533_/Q _1010_/Y _1014_/Y _1529_/Q _0996_/X _1015_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_34_241 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1292__A1 _1247_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1044__A1 _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1044__B2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1328__A1_N _0760_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1347__A2 _1339_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1490__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_333 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1551__D _1551_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_34 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_56 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0745__A usb_address[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1283__B2 _1240_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1035__A1 _0826_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1035__B2 _0840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1555__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1338__A2 _1337_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_63 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1461__D _1180_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_355 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_358 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1274__A1 _1420_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_200 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_233 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1026__B2 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1026__A1 _1020_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _1119_/Y _0920_/B rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1495_ _1495_/D _1495_/Q rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_119 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_141 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_185 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1546__D _1077_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_21 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1256__A1 _1245_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_391 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0922__B _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__B1 _1467_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_9 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1456__D _1456_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1192__B1 _1187_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1280_ _1423_/Q _1273_/X _0707_/C _1280_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_48_130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_339 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0832__B _0832_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0995_ _0823_/A _0823_/B _0992_/X _0993_/X _0994_/X _0995_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_8_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_292 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1004__A2_N _0840_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1547_ _1079_/X _1078_/A _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1478_ _1281_/X _0707_/D _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_39_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_358 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1238__B2 _1204_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1238__A1 _1603_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0742__B _1313_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_207 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1174__B1 _1581_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_314 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_317 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_125 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1570__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1229__A1 _1598_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0933__A _0869_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0988__B1 data_out[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_0780_ _0780_/A _1327_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_5_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_251 VGND VPWR sky130_fd_sc_hd__decap_3
X_1401_ _0887_/A _1399_/X _1401_/C _1401_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_1332_ _0771_/A _1340_/B _1330_/X _1331_/Y _1507_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__1551__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1263_ _1252_/B _1262_/X _1250_/C _1263_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0827__B _0827_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_122 VGND VPWR sky130_fd_sc_hd__fill_1
X_1194_ _1250_/C _1194_/B _1194_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_24_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0843__A _0843_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_350 VGND VPWR sky130_fd_sc_hd__fill_2
X_0978_ _0969_/X _0971_/X _1525_/Q _1440_/Q _0972_/X _0978_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_10_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_144 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_56 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0753__A _0734_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_309 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_361 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1424__CLK _1514_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0985__A3 _1444_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_99 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1574__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0928__A rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_239 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0735__A2_N _1447_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_158 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_383 VGND VPWR sky130_fd_sc_hd__fill_2
X_0901_ _0901_/A _0901_/B _1485_/Q _0901_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0813__D _1581_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0976__A3 _1523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0832_ _0821_/Y _0832_/B _0833_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1386__B1 _1388_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0763_ _0759_/X _0762_/X _0716_/X _0763_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_51_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1315_ _1315_/A _1315_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0897__C1 _0896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0838__A _1461_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0900__A3 _0786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_1246_ _0715_/B _1247_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1492__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1310__B1 _1309_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1177_ _0813_/C _1090_/X _1583_/Q _1092_/X _1177_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_109 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1447__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_136 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_180 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1597__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk_48 clkbuf_3_6_0_clk_48/X _1467_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1554__D _1554_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1509__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0748__A usb_address[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_283 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1301__B1 _1296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_32 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1298__B _0713_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_375 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1368__B1 _1363_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1464__D _1463_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1100_ _1557_/Q _1090_/X _0906_/A _1095_/X _1100_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_1031_ _0829_/X _0853_/A _0776_/B _0853_/Y _1031_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_46_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_106 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1071__A2 _1069_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1001__B _1056_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0815_ _0810_/X _0909_/C _0815_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1359__B1 _1355_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0746_ _0743_/Y _0744_/B _0745_/Y _1444_/Q _0746_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_217 VGND VPWR sky130_fd_sc_hd__fill_2
X_1229_ _1598_/Q _1216_/X _1228_/X _1229_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1399__A data_in[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1549__D _1549_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_172 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0750__B _0738_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_1_0_clk_48_A clkbuf_4_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1612__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0909__C _0909_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_261 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0925__B _0924_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_294 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1102__A _1102_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1459__D _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_297 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _1173_/X _0813_/A rst_n _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_14_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1014_ _1014_/A _1014_/B _1013_/X _0846_/C _1014_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__0835__B _0835_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1292__A2 tx_en VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1012__A _0818_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0851__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1044__A2 _0829_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0729_ _0755_/B _0895_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_57_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_267 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1035__A2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0761__A _0720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1533__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1596__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_146 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1524__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_220 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_264 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1274__A2 _1273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1508__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_256 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1026__A2 _0834_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1281__A2_N _1280_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1563_ _1563_/D _0919_/D rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1494_ _0796_/X _1357_/B rst_n _1514_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_39_345 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_326 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_59 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_clk_48 clkbuf_4_1_0_clk_48/A _1529_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_1_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1562__D _1562_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_67 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0756__A data_in_valid VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_197 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_318 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1256__A2 _1252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_245 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0922__C _0922_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_278 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0767__A1 _0766_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__B2 _0766_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1312__A1_N _1309_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1472__D _1192_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1192__A1 _0719_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_304 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_392 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1480__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0994_ _0994_/A _0994_/B _0994_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1404__C1 _1403_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_71 VGND VPWR sky130_fd_sc_hd__fill_2
X_1546_ _1077_/X _1002_/C _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1477_ _1279_/X _0707_/A _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_39_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_197 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_318 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1238__A2 _1204_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_392 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_329 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1200__A _1200_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0742__C _0739_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0749__A1 usb_address[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1557__D _1557_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_11 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1174__B2 _1092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1174__A1 _0813_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_18 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1229__A2 _1216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_370 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0933__B _1399_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0988__A1 _0901_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0988__B2 _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1110__A _1109_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1467__D rx_j VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_285 VGND VPWR sky130_fd_sc_hd__fill_2
X_1400_ _1425_/Q _1400_/B _1401_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_204 VGND VPWR sky130_fd_sc_hd__fill_2
X_1331_ _0771_/A _1340_/B _1331_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_1262_ _1250_/A _1245_/X _1262_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_1193_ _0873_/A _1250_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_36_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_104 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0843__B _0843_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_148 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1020__A _0823_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_395 VGND VPWR sky130_fd_sc_hd__fill_2
X_0977_ _0969_/X _0971_/X _1524_/Q _1439_/Q _0972_/X _1439_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_10_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_1529_ _1015_/X _1529_/Q rst_n _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_27_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0753__B _0753_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_218 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0928__B tx_en VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_148 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1083__B1 _1082_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0900_ _0785_/X _0889_/Y _0786_/Y _0891_/X _0899_/X _1488_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XPHY_90 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_170 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_0831_ _0829_/X _0830_/X _0829_/X _0830_/X _0843_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0762_ _0760_/Y _1185_/B _0762_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1386__A1 _1366_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1314_ _0958_/X _1313_/X _0935_/A _1503_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0897__B1 _0732_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_207 VGND VPWR sky130_fd_sc_hd__fill_2
X_1245_ _0874_/B _1245_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_49_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0842__A2_N _0841_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1176_ _1581_/Q _1171_/X _1175_/X _1582_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1310__A1 _0874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_284 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1310__B2 _1300_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_37 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0888__B1 _0887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0748__B _0747_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1570__D _1570_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_23 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1301__A1 _1259_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_67 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1541__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_354 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_314 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1368__B2 _1367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1368__A1 _0887_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0939__A _0938_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1480__D _1287_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1030_ _0835_/A _0853_/A _0776_/A _0853_/Y _1516_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_34_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0803__B1 _0798_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1001__C _1000_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0814_ _0811_/Y _0814_/B _0814_/C _0814_/D _0909_/C VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__1359__A1 _0886_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0745_ usb_address[1] _0745_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0849__A _1187_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1228_ _1228_/A _1222_/B _1228_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_26 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_262 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_284 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1564__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1159_ _1159_/A _0924_/X _1160_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1399__B _1399_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_243 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_287 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1047__B1 _1532_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1565__D _1122_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0734__A2_N _1443_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0759__A _0759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0909__D _0908_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1286__B1 _1285_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1038__B1 _1037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1475__D _1475_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1210__B1 _1207_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1437__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1587__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_251 VGND VPWR sky130_fd_sc_hd__fill_2
X_1013_ _0891_/X _1532_/Q _1013_/C _1013_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1277__B1 _0707_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_276 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1029__B1 _0840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0851__B _0816_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_93 VGND VPWR sky130_fd_sc_hd__decap_4
X_0728_ _0777_/A _0879_/A _0728_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_47 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1203__A _1202_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_246 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1564__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_98 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_397 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_276 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1026__A3 _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _1562_/D _0919_/C rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1493_ _1493_/D _1329_/A rst_n _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_39_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_335 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__B _0818_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_360 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_382 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0862__A _0862_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1602__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_79 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_390 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0772__A _0772_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_239 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0922__D _0922_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__A2 _0766_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1192__A2 _0718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0947__A endpoint[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_176 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_187 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_157 VGND VPWR sky130_fd_sc_hd__decap_4
X_0993_ _0891_/X _0846_/A _0818_/B _0993_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1404__B1 _1410_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1168__C1 _1167_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1486__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_1545_ _1075_/X _0999_/D _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1018__A _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1476_ _1277_/X _0707_/B _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0857__A _0816_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_341 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_227 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0742__D _0742_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__A2 _0747_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_36 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1573__D _1573_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1174__A2 _1090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_66 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_157 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0988__A2 _0970_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1110__B _1107_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_297 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1483__D _1312_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1330_ _1330_/A _1330_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_216 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_249 VGND VPWR sky130_fd_sc_hd__fill_2
X_1261_ _1258_/Y _1254_/X _1252_/A _1260_/Y _1261_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_1192_ _0719_/A _0718_/X _1187_/X _1192_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_24_308 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_371 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0843__C _0843_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_138 VGND VPWR sky130_fd_sc_hd__fill_2
X_0976_ _0969_/X _0971_/X _1523_/Q _1438_/Q _0972_/X _1438_/D VGND VPWR sky130_fd_sc_hd__a32o_4
X_1528_ _1019_/X _1528_/Q rst_n _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_238 VGND VPWR sky130_fd_sc_hd__fill_2
X_1459_ _1044_/X _0832_/B _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_27_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0753__C _0742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1568__D _1568_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1470__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1083__A1 _1003_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_341 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1478__D _1281_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0830_ _0823_/B _1037_/A _0830_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0761_ _0720_/X _1185_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1386__A2 _1382_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1313_ _1313_/A _0879_/A _1315_/A _1313_/D _1313_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0897__A1 _1316_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_219 VGND VPWR sky130_fd_sc_hd__fill_2
X_1244_ _1250_/A _1260_/B _0759_/X _1250_/C _1244_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1310__A2 _1245_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1175_ _0813_/C _1090_/A _1175_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_32_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_366 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0870__A data_in_valid VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_388 VGND VPWR sky130_fd_sc_hd__fill_1
X_0959_ _0855_/X _0955_/X _1435_/Q _1443_/Q _0958_/X _0959_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1493__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0888__A1 _1329_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1301__A2 _1300_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_127 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0964__A2_N _0962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1518__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0780__A _0780_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_388 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_326 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_29 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1368__A2 _1361_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1116__A _1128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0955__A _1413_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_288 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0803__B2 _0802_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A1 _0799_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1001__D _1001_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0813_ _0813_/A _0813_/B _0813_/C _1581_/Q _0814_/D VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1359__A2 _1354_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0744_ _0743_/Y _0744_/B _0744_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1227_ _1597_/Q _1216_/X _1226_/X _1227_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_1158_ _1158_/A _1155_/Y _1158_/C _1575_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_25_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_266 VGND VPWR sky130_fd_sc_hd__fill_2
X_1089_ _1016_/X _1088_/X _1552_/Q _1016_/X _1552_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_299 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1611__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1047__B2 _1046_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_185 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1581__D _1174_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_45 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0775__A _0774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1286__A1 _1284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_200 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_255 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1038__A1 _1036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_134 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_81 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1210__B2 _1204_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1210__A1 _1207_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1491__D _1491_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_358 VGND VPWR sky130_fd_sc_hd__decap_8
X_1012_ _0818_/B _1014_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1277__B2 _1241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_266 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1029__A1 _1527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1029__B2 _1021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0851__C _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VPWR sky130_fd_sc_hd__decap_4
X_0727_ _1492_/Q _0879_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0960__B1 _1444_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1531__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_299 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1576__D _1163_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_303 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_91 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1486__D _0915_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1561_ _1108_/X _0919_/B rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1554__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_1492_ _1492_/D _1492_/Q rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_39_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_358 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__C _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_391 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1049__A1_N _1048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1214__A _1593_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_203 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0772__B _0772_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1427__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1577__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1177__B1 _1583_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0947__B _0945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1101__B1 _0907_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0992_ _0994_/B _0992_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_44_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1404__A1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1168__B1 _1147_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1544_ _1073_/X _1072_/A _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_5_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0915__B1 _1484_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1475_ _1475_/D _1269_/A _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_39_111 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1034__A _1014_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0873__A _0873_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_191 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_7 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0783__A _1327_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_342 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0988__A3 _1447_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1398__B1 _1424_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1119__A _1128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0958__A _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1260_ _1259_/X _1260_/B _1260_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_1191_ _0719_/A _1189_/Y _1190_/X _1187_/X _1191_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_36_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_320 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0843__D _0842_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0975_ _0969_/X _0971_/X _1522_/Q _1437_/Q _0972_/X _0975_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_1527_ _1527_/D _1527_/Q rst_n _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__0868__A _0724_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1458_ _1458_/D _0829_/B _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_67_283 VGND VPWR sky130_fd_sc_hd__decap_4
X_1389_ handshake[1] _0720_/X _0759_/X _1389_/D _1389_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_27_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0753__D _0753_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_183 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1584__D _1178_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_268 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0778__A _1358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1304__B1 _0712_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1539__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1083__A2 _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_81 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_92 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1121__B1_N _1120_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0760_ handshake[1] _0760_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1494__D _0796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_91 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0897__A2 _0895_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1312_ _1309_/Y _1296_/X _1296_/X tx_j _1312_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_41 VGND VPWR sky130_fd_sc_hd__fill_2
X_1243_ _0874_/C _0715_/B _1260_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_49_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_231 VGND VPWR sky130_fd_sc_hd__decap_4
X_1174_ _0813_/A _1090_/X _1581_/Q _1092_/X _1174_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_64_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_323 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_356 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0870__B _0887_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0958_ _0957_/X _0958_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0889_ _0789_/X _0889_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0888__A2 _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_117 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1222__A _1596_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_13 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1579__D _1170_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_378 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_338 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1368__A3 _1363_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1558__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1116__B _1115_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_401 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1132__A _1131_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_245 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1489__D _0765_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0971__A _0970_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A2 _0800_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0812_ _1583_/Q _0814_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_52_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_0743_ usb_address[5] _0743_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_1226_ _1598_/Q _1222_/B _1226_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1157_ _1155_/A _1156_/Y _1155_/B _1158_/C VGND VPWR sky130_fd_sc_hd__o21a_4
X_1088_ _1086_/Y _1059_/Y _1086_/A _1004_/X _1088_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0881__A _1358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1460__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_164 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1217__A _1217_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1286__A2 _1247_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_234 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1038__A2 _0827_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0791__A _0791_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_278 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_120 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1210__A2 _1204_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_1011_ _1534_/Q _1014_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_19_275 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_297 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1483__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_245 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_256 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1029__A2 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0851__D _0851_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_73 VGND VPWR sky130_fd_sc_hd__decap_3
X_0726_ _1317_/A _0755_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0960__B2 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0960__A1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0963__A2_N _0962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1037__A _1037_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0876__A _1187_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1209_ _1207_/Y _1208_/X _1589_/Q _1208_/X _1590_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_245 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1279__A1_N _1272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1592__D _1213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_78 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_67 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_366 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0786__A _0722_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_381 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1573__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_237 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1410__A _1350_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1502__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ _1104_/Y _1560_/Q rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_3_160 VGND VPWR sky130_fd_sc_hd__fill_2
X_1491_ _1491_/D _1319_/A rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_66_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_307 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__D _0846_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0_0_clk_48_A clkbuf_4_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_237 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_248 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_29 VGND VPWR sky130_fd_sc_hd__decap_4
X_0709_ _1606_/Q _1605_/Q _0709_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_1_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1214__B _1214_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_156 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0772__C _0772_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1230__A _1600_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1587__D _1184_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_281 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1177__B2 _1092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1177__A1 _0813_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_115 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1101__B2 _1092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_373 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1101__A1 _0906_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0991_ _0901_/A _0970_/X _1450_/Q data_out[7] _0961_/X _1434_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1497__D _1497_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0860__B1 _1413_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1404__A2 _1402_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_292 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1521__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_1612_ _1612_/D _1612_/Q rst_n _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1168__A1 _0916_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_52 VGND VPWR sky130_fd_sc_hd__decap_4
X_1543_ _1071_/X _0999_/B _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1474_ _1271_/X _1201_/A _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0915__B2 _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_123 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1315__A _1315_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_167 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_318 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_340 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1495__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_35 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_318 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0783__B _0783_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1544__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_310 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0842__B1 _0837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1398__A1 _0887_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1398__B2 _1397_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1119__B _1119_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_60 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_218 VGND VPWR sky130_fd_sc_hd__decap_12
X_1190_ _0717_/A _1186_/A _1190_/X VGND VPWR sky130_fd_sc_hd__and2_4
Xclkbuf_3_1_0_clk_48 clkbuf_3_1_0_clk_48/A clkbuf_4_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_17_340 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_181 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_354 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_398 VGND VPWR sky130_fd_sc_hd__fill_2
X_0974_ _0969_/X _0971_/X _1521_/Q _1436_/Q _0972_/X _0974_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_1526_ _1028_/X _1526_/Q rst_n _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1457_ _1042_/X _0825_/B _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1388_ _1388_/A _1388_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1605__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1567__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_159 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1077__B1 _1076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_170 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_343 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0778__B _0778_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_240 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_115 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1304__A1 _1305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0794__A _1313_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1068__B1 _1067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_321 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_195 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0969__A _1187_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1311_ _1309_/Y _1300_/X _1310_/X tx_j VGND VPWR sky130_fd_sc_hd__a21bo_4
X_1242_ _0874_/B _1252_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_2_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_273 VGND VPWR sky130_fd_sc_hd__decap_3
X_1173_ _0813_/B _1171_/X _1172_/X _1173_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_64_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0870__C _0870_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0957_ _0891_/X _0957_/B _0957_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1231__B1 _1230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_0888_ _1329_/A _0876_/X _0887_/X _1493_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0879__A _0879_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1545__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1509_ _1509_/D _1509_/Q rst_n _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_28_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_405 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1222__B _1222_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1595__D _1221_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0789__A _0788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1527__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1413__A _0856_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_298 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_0811_ _0811_/A _0811_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1213__B1 _1212_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0742_ _0736_/Y _1313_/A _0739_/X _0742_/D _0742_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_6_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1225_ _1596_/Q _1216_/X _1224_/X _1225_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_1156_ _0917_/X _1156_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_37_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1307__A2_N _1306_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1087_ _1086_/Y _1057_/X _1550_/Q _1057_/X _1551_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1605__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0881__B _0881_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_154 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_4_0_clk_48 clkbuf_4_5_0_clk_48/A _1583_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1217__B _1214_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_243 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_276 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1408__A _1289_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1591__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_349 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1143__A _1143_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1010_ _1009_/X _1010_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0725_ _0716_/X _0725_/B _0886_/A _0725_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_6_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1318__A _1318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0960__A2 _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1037__B _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0876__B tx_en VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_338 VGND VPWR sky130_fd_sc_hd__fill_2
X_1208_ _1205_/A _1208_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_360 VGND VPWR sky130_fd_sc_hd__fill_2
X_1139_ _0925_/Y _1138_/X _1139_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0892__A _0892_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_268 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1228__A _1228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_323 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1601__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_50 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_216 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1416__B1 _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1410__B _1410_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_71 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1138__A _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_172 VGND VPWR sky130_fd_sc_hd__decap_3
X_1490_ _0878_/X _0892_/A rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1450__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_146 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_363 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1407__B1 data_in[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_293 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1048__A _1533_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0708_ _1285_/A _0708_/B _1482_/Q _0708_/D _0715_/B VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1170__A2_N _0841_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0887__A _0887_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_113 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1343__C1 _1342_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_37 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0772__D _1512_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1230__B _1222_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_249 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1177__A2 _1090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0797__A _1463_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1473__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1334__C1 _1333_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_382 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1101__A2 _1090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_396 VGND VPWR sky130_fd_sc_hd__fill_1
X_0990_ _0901_/A _0970_/X _1449_/Q data_out[6] _0961_/X _0990_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__0860__A1 _0732_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_81 VGND VPWR sky130_fd_sc_hd__decap_3
X_1611_ _1306_/Y _0712_/B rst_n _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1168__A2 _1166_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1542_ _1068_/X _0999_/C _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_5_75 VGND VPWR sky130_fd_sc_hd__fill_2
X_1473_ _1473_/D _1473_/Q _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_54_127 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0915__A2_N _0913_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1331__A _0771_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_396 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1496__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_127 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1241__A _1240_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_363 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1598__D _1227_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_193 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_322 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0842__B2 _0841_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_399 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1398__A2 _0758_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_374 VGND VPWR sky130_fd_sc_hd__fill_2
X_0973_ _0969_/X _0971_/X _1520_/Q _1435_/Q _0972_/X _1435_/D VGND VPWR sky130_fd_sc_hd__a32o_4
X_1525_ _1525_/D _1525_/Q rst_n _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_19_29 VGND VPWR sky130_fd_sc_hd__decap_3
X_1456_ _1456_/D _0836_/B _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1387_ data_in[3] _1399_/B _1387_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1077__A1 _0999_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_311 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_38 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1236__A _1603_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1511__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1304__A2 _1296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0794__B _0794_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1068__A1 _1001_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_333 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_174 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0751__B1 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_270 VGND VPWR sky130_fd_sc_hd__fill_2
X_1310_ _0874_/A _1245_/X _1309_/Y _1300_/X _1310_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_1_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_32 VGND VPWR sky130_fd_sc_hd__fill_2
X_1241_ _1240_/X _1241_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1172_ _0813_/A _1090_/A _1172_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_66_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_296 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_244 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_369 VGND VPWR sky130_fd_sc_hd__fill_2
X_0956_ _1413_/B _0957_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1231__A1 _1228_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0887_ _0887_/A _0887_/B _0756_/Y _0887_/D _0887_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0990__B1 data_out[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0879__B _0879_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1056__A _1056_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1534__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1508_ _1334_/X _0771_/B rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1439_ _1439_/D _1439_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0895__A _1317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_41 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0746__A2_N _0744_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1047__A1_N _1046_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1567__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1413__B _1413_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_225 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1551__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0810_ _1587_/Q _1183_/B _0810_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1213__A1 _1591_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0741_ usb_address[3] _0740_/Y usb_address[3] _0740_/Y _0742_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1557__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_1224_ _1597_/Q _1222_/B _1224_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1155_ _1155_/A _1155_/B _1155_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_1086_ _1086_/A _1086_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_16_19 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_277 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0881__C _0864_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_0939_ _0938_/X _0945_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0963__B1 _1437_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1140__B1 _1158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_225 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0954__B1 _0953_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1408__B _1381_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_211 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1143__B _1139_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_280 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1198__B1 _1252_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0724_ _0724_/A _0886_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0960__A3 _1436_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1489__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_1207_ _1207_/A _1207_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_27_29 VGND VPWR sky130_fd_sc_hd__decap_3
X_1138_ _0922_/A _0922_/B _0922_/D _0918_/B _1138_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0892__B _0892_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1069_ _0994_/B _1069_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_43_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_291 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0936__B1 _0935_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1228__B _1222_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_335 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_350 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1113__B1 _1158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_95 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1416__A1 _1414_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_50 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1138__B _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1582__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1154__A _1154_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1511__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1352__B1 _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_317 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_386 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1407__A1 _1389_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1407__B2 _0758_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1329__A _1329_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0707_ _0707_/A _0707_/B _0707_/C _0707_/D _0708_/D VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0887__B _0887_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1064__A _0818_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1343__B1 _1330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_16 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1334__B1 _1330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_331 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0860__A2 _0856_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_243 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1149__A _1148_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_1610_ _1303_/X _1305_/A rst_n _1611_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1541_ _1541_/D _1001_/D _0927_/X _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1472_ _1192_/X _0719_/A _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1325__B1 _1324_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_331 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1331__B _1340_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_389 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1059__A _1004_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0898__A _1492_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1398__A3 data_in[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_213 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1440__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1590__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1307__B1 _1612_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_334 VGND VPWR sky130_fd_sc_hd__fill_2
X_0972_ _0961_/X _0972_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1524_ _1026_/X _1524_/Q rst_n _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1455_ _1040_/X _0834_/B _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_67_242 VGND VPWR sky130_fd_sc_hd__fill_2
X_1386_ _1366_/X _1382_/X _1388_/A _1386_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1342__A _1342_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_29 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1077__A2 _1069_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_150 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1463__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_131 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_7 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_238 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0794__C _0728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1252__A _1252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1068__A2 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1277__A1_N _1272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_142 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_9 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0751__A1 _0745_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_22 VGND VPWR sky130_fd_sc_hd__fill_1
X_1240_ _0715_/C _1240_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_49_242 VGND VPWR sky130_fd_sc_hd__fill_2
X_1171_ _1092_/X _1171_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_64_223 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1162__A _1159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1486__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_186 VGND VPWR sky130_fd_sc_hd__fill_2
X_0955_ _1413_/B _0955_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1231__A2 _1205_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0886_ _0886_/A _0887_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0990__A1 _0901_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0990__B2 _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1507_ _1507_/D _0771_/A rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1061__A2_N _1060_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1438_ _1438_/D _1438_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0895__B _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1072__A _1072_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1369_ _0758_/Y _1362_/X _1369_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_197 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1247__A _0874_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1213__A2 _1208_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0740_ _1446_/Q _0740_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_6_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_1223_ _1595_/Q _1216_/X _1222_/X _1596_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_28_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_223 VGND VPWR sky130_fd_sc_hd__decap_4
X_1154_ _1154_/A _1154_/B _1155_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_37_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_1085_ _1002_/D _1039_/X _1084_/X _1550_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_52_248 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_270 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_101 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_189 VGND VPWR sky130_fd_sc_hd__decap_4
X_0938_ _0937_/X _0938_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1501__CLK _1514_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0963__B2 _0962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1067__A _0999_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0869_ _0869_/A _0716_/X _0870_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1140__A1 _1137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_259 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_112 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_270 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_138 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0954__A1 _1437_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_248 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1524__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_87 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1198__A1 _1473_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0723_ _0722_/X _0725_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_1206_ _1214_/B _1204_/Y _1589_/Q _1205_/X _1589_/D VGND VPWR sky130_fd_sc_hd__o22a_4
X_1137_ _1137_/A _1137_/B _1137_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_25_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1350__A _1495_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1068_ _1001_/D _1057_/X _1067_/X _1068_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1500__D _0954_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_270 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0936__A1 _1506_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1113__A1 _1110_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1547__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_226 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1260__A _1259_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1416__A2 _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_229 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1138__C _0922_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1352__A1 _1350_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1154__B _1154_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1352__B2 _1185_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_321 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1407__A2 _1406_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_240 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1329__B _1329_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1040__B1 _0834_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0706_ _0759_/A _0715_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0887__C _0756_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1343__A1 _0772_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_332 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1080__A _1003_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_354 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0854__B1 _0853_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1031__B1 _0776_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1334__A1 _0771_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_192 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1098__B1 _1556_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1149__B _1149_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_1540_ _1540_/D _1540_/Q _0927_/X _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1022__B1 _1520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1165__A _1164_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1471_ _1191_/X _0717_/A _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1325__A1 _0867_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1089__B1 _1552_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_310 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_313 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1261__B1 _1252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0898__B _0898_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_27 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_181 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_335 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_346 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_64 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1004__B1 _1552_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1307__B2 _1306_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_346 VGND VPWR sky130_fd_sc_hd__fill_2
X_0971_ _0970_/X _0971_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1534__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_390 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1597__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0999__A _1540_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1523_ _1523_/D _1523_/Q rst_n _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1454_ _1038_/X _1037_/A _1454_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_4_280 VGND VPWR sky130_fd_sc_hd__fill_2
X_1385_ _1421_/Q _1397_/B _1383_/X _1384_/X _1385_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_27_107 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1608__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_265 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0794__D _1313_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1252__B _1252_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1244__A2_N _1260_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_63 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_85 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_96 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1225__B1 _1224_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_95 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0751__A2 _1444_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_45 VGND VPWR sky130_fd_sc_hd__decap_4
X_1170_ _1094_/X _0841_/Y _0813_/B _1094_/X _1170_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1162__B _0924_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_327 VGND VPWR sky130_fd_sc_hd__fill_1
X_0954_ _1437_/Q _0942_/X _0953_/X _0954_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0885_ _0885_/A _0884_/Y _1491_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0990__A2 _0970_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1506_ _1506_/D _1506_/Q rst_n _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1437_ _0975_/X _1437_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0895__C _0754_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1368_ _0887_/A _1361_/X _1363_/X _1363_/A _1367_/X _1368_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_55_213 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1072__B _1064_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1430__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_235 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1503__D _1503_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1299_ _1201_/A _1196_/Y _1604_/Q _1196_/Y _1299_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1580__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_132 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_338 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_clk_48 clkbuf_2_1_0_clk_48/A clkbuf_3_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1247__B _0874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1576__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_320 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1505__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1453__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1222_ _1596_/Q _1222_/B _1222_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1153_ _1154_/A _1154_/B _1147_/A _1152_/Y _1153_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_1084_ _1550_/Q _1014_/B _1084_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_60_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_146 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_168 VGND VPWR sky130_fd_sc_hd__decap_4
X_0937_ _0891_/X _1492_/Q _1313_/D _0937_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__1067__B _1064_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0868_ _0724_/A _0869_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0799_ _1466_/Q _0799_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_28_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1140__A2 _1139_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_249 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_260 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1258__A _1329_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0954__A2 _0942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1476__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_371 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_393 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_279 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_71 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1198__A2 _1196_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0722_ _0721_/X _0722_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0800__A _1466_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1205_ _1205_/A _1205_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1136_ _0918_/B _1137_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_25_205 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_249 VGND VPWR sky130_fd_sc_hd__fill_1
X_1067_ _0999_/C _1064_/X _1067_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1498__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1078__A _1078_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1499__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0936__A2 _0870_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0710__A _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_304 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_308 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1113__A2 _1111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1260__B _1260_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_271 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1138__D _0918_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_164 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1352__A2 _1351_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_71 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_7 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4_0_clk_48 clkbuf_3_5_0_clk_48/A clkbuf_4_9_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1601__D _1233_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_377 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1520__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1407__A3 _1399_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1040__B2 _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1040__A1 _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0887__D _0887_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1343__A2 _0772_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1484__SET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1361__A data_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1080__B _1014_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1608__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_1119_ _1128_/A _1119_/B _1119_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__1511__D _1345_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0854__A1 _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_296 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1031__A1 _0829_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1031__B2 _0853_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0790__B1 _0786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1514__CLK _1514_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1334__A2 _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_63 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1098__A1 _1555_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_322 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1098__B2 _1095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1421__D _1385_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_201 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_296 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_234 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1022__B2 _1021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1022__A1 _1020_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_89 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_56 VGND VPWR sky130_fd_sc_hd__fill_1
X_1470_ _1470_/D _1470_/Q _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_67_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1325__A2 _1321_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1181__A _1588_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1089__B2 _1016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_322 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_171 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1261__B2 _1260_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1261__A1 _1258_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1537__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1506__D _1506_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1599_ _1229_/X _1228_/A _0928_/X _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1091__A _1090_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_311 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_21 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1004__B2 _0840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1266__A _1265_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0763__B1 _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_163 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_399 VGND VPWR sky130_fd_sc_hd__fill_2
X_0970_ _1413_/B _0970_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0999__B _0999_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1522_ _1024_/X _1522_/Q rst_n _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1453_ _1035_/X _0826_/B _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1384_ data_in[2] _0935_/Y _1384_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_196 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_144 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0993__B1 _0818_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1086__A _1086_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_clk_48 clkbuf_4_7_0_clk_48/A _1575_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_200 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1170__B1 _0813_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_288 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1540__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_20 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_325 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_100 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1225__A1 _1596_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0984__B1 data_out[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_152 VGND VPWR sky130_fd_sc_hd__fill_2
X_0953_ endpoint[3] _0945_/B _0953_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0975__B1 _1437_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0884_ _1329_/A _0892_/B _1319_/A _0775_/X _0884_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XANTENNA__0990__A3 _1449_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1505_ _1353_/X _0759_/A rst_n _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1436_ _0974_/X _1436_/Q _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1367_ _1364_/X _1366_/X _1367_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_258 VGND VPWR sky130_fd_sc_hd__fill_2
X_1298_ _0712_/A _0713_/A _1298_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_23_100 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0966__B1 _0744_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0713__A _0713_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1247__C _1245_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_73 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1221_ _1217_/A _1216_/X _1220_/X _1221_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1604__D _1239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_203 VGND VPWR sky130_fd_sc_hd__fill_2
X_1152_ _1154_/A _1150_/X _1152_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_37_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_206 VGND VPWR sky130_fd_sc_hd__fill_2
X_1083_ _1003_/A _1039_/X _1082_/X _1549_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_37_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_291 VGND VPWR sky130_fd_sc_hd__fill_2
X_0936_ _1506_/Q _0870_/C _0935_/Y _1506_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_9_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0948__B1 _0947_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0867_ _0760_/Y _0867_/B _0887_/D VGND VPWR sky130_fd_sc_hd__and2_4
X_0798_ _0798_/A _0798_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_1419_ _1368_/X _1363_/A _1514_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1514__D _1325_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_247 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0708__A _1285_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_269 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_103 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_283 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_107 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1364__B1 _1357_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_350 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1424__D _1424_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_250 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_283 VGND VPWR sky130_fd_sc_hd__fill_2
X_0721_ _0759_/A _0720_/X _0721_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1420__CLK _1514_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1570__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1204_ _1204_/A _1204_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_65_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_1135_ _0922_/B _1131_/X _1147_/A _1137_/B _1135_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_1066_ _1540_/Q _1057_/X _1065_/X _1541_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_18_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1078__B _1014_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1509__D _1509_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0919_ _1560_/Q _0919_/B _0919_/C _0919_/D _0920_/C VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1094__A _1090_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_191 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_87 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_20 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1443__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1269__A _1269_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1419__D _1368_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1593__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0901__A _0901_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1337__B1 _0772_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_356 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_294 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1275__A1_N _1272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1560__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1040__A2 _0830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0811__A _0811_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1328__B1 _1315_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_331 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1361__B _1399_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_386 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1466__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1118_ _0920_/B _1114_/X _1117_/X _1119_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XANTENNA__0854__A2 _0818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_209 VGND VPWR sky130_fd_sc_hd__fill_2
X_1049_ _1048_/Y _1036_/X _1532_/Q _1036_/X _1533_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_253 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0721__A _0759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1031__A2 _0853_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0790__B2 _0789_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_109 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_353 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_386 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1098__A2 _1094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_356 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_378 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1089__A2_N _1088_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_84 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1022__A2 _0832_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1489__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1181__B _1187_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1612__D _1612_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_131 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0806__A _0806_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1261__A2 _1254_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1598_ _1227_/X _1598_/Q _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1522__D _1024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_164 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_367 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0716__A _0757_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_98 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0763__A1 _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_41 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1432__D _0989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_131 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_186 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0999__C _0999_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1521_ _1521_/D _1521_/Q rst_n _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1607__D _1607_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1452_ _1415_/X _0856_/B _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1383_ _1421_/Q _1409_/B _1382_/X _1383_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_67_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_315 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_348 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1504__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0790__A2_N _0786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1367__A _1364_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A1 _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_208 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1517__D _1031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_109 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1170__B2 _1094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_21 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_112 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_87 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1225__A2 _1216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_370 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0984__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0984__B2 _0981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1427__D _1427_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_61 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1527__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_123 VGND VPWR sky130_fd_sc_hd__fill_2
X_0952_ _1436_/Q _0942_/X _0951_/X _0952_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_20_318 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_330 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0975__B2 _0972_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0975__A1 _0969_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0883_ tx_en _0892_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1187__A _1187_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1504_ _1504_/D success rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1435_ _1435_/D _1435_/Q _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1366_ _1350_/X _0725_/B _1410_/B _1366_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_1297_ _1305_/A _1296_/X _1303_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_63_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_318 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0966__A1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0713__B _1300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0966__B2 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1247__D _1247_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1411__A2_N _0725_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_259 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_229 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_145 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0904__A _0904_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1585__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_1220_ _1595_/Q _1222_/B _1220_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1514__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_1151_ _1149_/X _1150_/X _1158_/A _1573_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1082_ _1002_/D _1014_/B _1082_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_60_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0814__A _0811_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0935_ _0935_/A _0935_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0948__A1 _1450_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_171 VGND VPWR sky130_fd_sc_hd__fill_2
X_0866_ handshake[0] _0867_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_0797_ _1463_/Q _0797_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_1418_ _1605_/Q _1605_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_68_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_1349_ _1513_/Q _0773_/X _1330_/X _1513_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_28_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1380__A _1380_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__B _0708_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0884__B1 _1319_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1530__D _1530_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_270 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_clk_48_A clkbuf_3_7_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0724__A _0724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_11 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1061__B1 _1539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1364__A1 _0725_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1290__A _1289_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1440__D _0978_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_13 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1052__B1 _1051_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0720_ _0719_/X _0720_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_10_181 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1203_ _1202_/X _1204_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_310 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0809__A _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_343 VGND VPWR sky130_fd_sc_hd__fill_2
X_1134_ _0922_/A _0922_/B _0922_/D _1150_/B _1137_/B VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_65_376 VGND VPWR sky130_fd_sc_hd__decap_12
X_1065_ _1001_/D _1064_/X _1065_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_21_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1291__B1 _1285_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1043__B1 _0829_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0918_ _0918_/A _0918_/B _0922_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1375__A _1409_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0849_ _1187_/A _0901_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1525__D _1525_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_332 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0719__A _0719_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_33 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_99 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1282__B1 _0708_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_406 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1269__B _1269_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_54 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_100 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1285__A _1285_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0901__B _0901_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1337__A1 _1335_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1435__D _1435_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_262 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1025__B1 _1523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_276 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1195__A _1194_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1328__B2 _1327_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_173 VGND VPWR sky130_fd_sc_hd__fill_2
X_1117_ _0920_/B _0920_/C _0925_/Y _1117_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_38_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91 VGND VPWR sky130_fd_sc_hd__fill_2
X_1048_ _1533_/Q _1048_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1264__B1 _1263_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0721__B _0720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_376 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1255__B1 _1254_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_64 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_75 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1560__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_247 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0912__A _0818_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1022__A3 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1191__C1 _1187_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0806__B _0805_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0822__A _0821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1597_ _1225_/X _1597_/Q _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1433__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1583__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1237__B1 _1234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__C1 _0993_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0732__A _0732_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0763__A2 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0907__A _1555_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0911__A2_N _0901_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_382 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0999__D _0999_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1520_ _1022_/X _1520_/Q rst_n _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1456__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1451_ _1451_/D _1414_/A _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1382_ _1357_/B _1381_/X _1382_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_67_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_279 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0817__A _0816_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1367__B _1366_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A2 _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1533__D _1533_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0727__A _1492_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_22 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_33 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_187 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_55 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_77 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_66 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0984__A2 _0980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1479__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_231 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_264 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1443__D _0959_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_110 VGND VPWR sky130_fd_sc_hd__fill_2
X_0951_ endpoint[2] _0945_/B _0951_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_13_371 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0975__A2 _0971_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0882_ _0879_/Y _0881_/X _0885_/A _1492_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_40_190 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1187__B _1187_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1385__C1 _1384_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1503_ _1503_/D data_strobe rst_n _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_4_9_0_clk_48_A clkbuf_4_9_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1434_ _1434_/D data_out[7] _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1365_ _0869_/A _0872_/X _1410_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_1296_ _1305_/B _1296_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_63_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_168 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0966__A2 _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1528__D _1019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1288__A _1482_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0904__B _0904_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1438__D _1438_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0920__A _0920_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_7 VGND VPWR sky130_fd_sc_hd__decap_3
X_1150_ _1154_/B _1150_/B _1150_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_1081_ _1078_/A _1069_/X _1080_/X _1081_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1554__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0814__B _0814_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0934_ _0933_/X _0935_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0948__A2 _0942_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0865_ _1492_/Q _0879_/B _1319_/A _0864_/Y _0865_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0830__A _0823_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0796_ _0785_/X _0790_/X _0794_/Y _0795_/X _0796_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_1417_ _1606_/Q _1605_/Q _1296_/X _1417_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_68_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_1348_ _1513_/Q _1346_/Y _1347_/X _1330_/X _1512_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0708__C _1482_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1279_ _1272_/X _1278_/Y _0707_/A _1240_/X _1279_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__0884__B2 _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0884__A1 _1329_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1058__A1_N _1056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_282 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1061__B2 _1016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_45 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_56 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0740__A _1446_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1517__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1364__A2 _0889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1290__B _1247_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_15_0_clk_48_A clkbuf_3_7_0_clk_48/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_296 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1052__A1 _1046_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1202_ _1196_/Y _1202_/B _1202_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_19_3 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_clk_48 clkbuf_0_clk_48/X clkbuf_2_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1133_ _0922_/A _1130_/B _1147_/A _1132_/Y _1568_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_65_388 VGND VPWR sky130_fd_sc_hd__decap_12
X_1064_ _0818_/B _1064_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0825__A _0821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1291__A1 _1288_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1291__B2 _1241_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0917_ _0916_/X _0917_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1043__B2 _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1043__A1 _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1375__B _1372_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0848_ _0777_/A _1187_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0779_ _0779_/A _0780_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1391__A _0758_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_182 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_322 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0719__B _0718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1541__D _1541_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_377 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_263 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1282__A1 _1424_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_285 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0901__C _1485_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1546__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_134 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1337__A2 _1336_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_171 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1451__D _1451_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_244 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1025__A1 _1020_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1025__B2 _1021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0784__B1 _0783_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_1116_ _1128_/A _1115_/Y _1563_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_53_336 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_358 VGND VPWR sky130_fd_sc_hd__fill_2
X_1047_ _1046_/X _1010_/Y _1532_/Q _1046_/X _1532_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_211 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1264__A1 _1241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1536__D _1054_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1255__A1 _1252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_204 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1007__A1 _0791_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1296__A _1305_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1446__D _0964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1191__B1 _1190_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_7 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_122 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_336 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_358 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_177 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_317 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_328 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_281 VGND VPWR sky130_fd_sc_hd__fill_2
X_1596_ _1596_/D _1596_/Q _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1592__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_185 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_339 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1237__B2 _1208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__B1 _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0732__B _0776_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_207 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1491__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1173__B1 _1172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_336 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0907__B _0905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_358 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_12_0_clk_48 clkbuf_3_6_0_clk_48/X _1577_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_380 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0923__A _1573_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__B1 data_out[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_361 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_394 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1579__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1508__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1209__A2_N _1208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_1450_ _0968_/X _1450_/Q _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1602__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1381_ _1381_/A _0722_/X _1381_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0911__B1 _1484_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0978__B1 _1440_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0833__A _0833_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_350 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_372 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_203 VGND VPWR sky130_fd_sc_hd__fill_2
X_1579_ _1170_/X _0813_/B rst_n _1583_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1550__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_291 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0743__A usb_address[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_11 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0984__A3 _1443_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1180__A2_N _1171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1146__B1 _1145_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_49 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0918__A _0918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_310 VGND VPWR sky130_fd_sc_hd__fill_2
X_0950_ _1435_/Q _0942_/X _0949_/X _1498_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1423__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0975__A3 _1522_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0881_ _1358_/A _0881_/B _0864_/B _0881_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__1187__C _1187_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1385__B1 _1383_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1573__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1502_ _0944_/Y setup rst_n _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1433_ _0990_/X data_out[6] _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_49_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1364_ _0725_/B _0889_/Y _1357_/B _1364_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_1295_ _0713_/A _1305_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_239 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0966__A3 _1440_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1376__B1 _1374_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1394__A _1350_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_9 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1544__D _1073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0738__A _1445_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1446__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_87 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1596__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0920__B _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1454__D _1038_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0878__C1 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1080_ _1003_/A _1014_/B _1080_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_33_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_220 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_clk_48 clkbuf_3_7_0_clk_48/A clkbuf_3_7_0_clk_48/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_60_242 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1523__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0814__C _0814_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0933_ _0869_/A _1399_/B _0933_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1087__A2_N _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0864_ _0861_/Y _0864_/B _0864_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0830__B _1037_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0795_ _0715_/A _1185_/B _0724_/A handshake[1] _0795_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_1416_ _1414_/A _0955_/X _0885_/A _1451_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_68_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_1347_ _0772_/C _1339_/X _1512_/Q _1347_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_68_397 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_228 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1469__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1278_ _1388_/A _1273_/X _0707_/D _1278_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__0884__A2 _0892_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__D _0708_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1389__A handshake[1] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_264 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1539__D _1539_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1349__B1 _1330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_397 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_261 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_clk_48 clkbuf_4_1_0_clk_48/A _1454_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1449__D _0967_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1052__A2 _1050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0931__A _0874_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1103__A1_N _1560_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1201_ _1201_/A _1604_/Q _1202_/B VGND VPWR sky130_fd_sc_hd__xnor2_4
XANTENNA__1611__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_356 VGND VPWR sky130_fd_sc_hd__fill_2
X_1132_ _1131_/X _1132_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_65_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_1063_ _1539_/Q _1057_/X _1062_/X _1540_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_18_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0825__B _0825_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1002__A _1072_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1291__A2 _1267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0916_ _0916_/A _1159_/A _0916_/C _0916_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1043__A2 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0841__A _0840_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0847_ _1485_/Q _0818_/X _0846_/X _0847_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__1375__C _0935_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0778_ _1358_/A _0778_/B _0779_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1391__B _1391_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_209 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1282__A2 _1273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_312 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0926__A _0925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_337 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0741__A2_N _0740_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1025__A2 _0836_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0784__A1 _0769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_109 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_312 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_142 VGND VPWR sky130_fd_sc_hd__fill_2
X_1115_ _0919_/D _1111_/X _1114_/X _1115_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XANTENNA__0836__A _0821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1046_ _0912_/X _1046_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1507__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_201 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1264__A2 _1261_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1552__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1552__D _1552_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1255__A2 _1196_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_65 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_238 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1007__A2 _0996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1412__C1 _1411_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_38 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1191__A1 _0719_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1462__D rx_se0 VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_293 VGND VPWR sky130_fd_sc_hd__fill_2
X_1595_ _1221_/X _1595_/Q _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_26_315 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_348 VGND VPWR sky130_fd_sc_hd__fill_2
X_1029_ _1527_/Q _1018_/X _0840_/X _1021_/X _1527_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_41_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_58 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1397__A _1364_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__A1 _0901_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1547__D _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1173__A1 _0813_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0907__C _0906_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_167 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0923__B _1145_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__B2 _0981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1457__D _1042_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_252 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_1380_ _1380_/A _1409_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_67_237 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0911__B2 _0910_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_148 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0978__A1 _0969_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0978__B2 _0972_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1010__A _1009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_1578_ _1578_/D _0916_/C rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_66_270 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_24 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_329 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_35 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_57 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_57 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_362 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1146__A1 _1145_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_207 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0918__B _0918_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_292 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_156 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0934__A _0933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_340 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_362 VGND VPWR sky130_fd_sc_hd__decap_4
X_0880_ _0880_/A _0783_/B _0881_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1385__A1 _1421_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1501_ _0946_/X direction_in rst_n _1514_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1432_ _0989_/X data_out[5] _1443_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1363_ _1363_/A _1362_/X _0758_/Y _1363_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__0896__B1 _0776_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1294_ _1506_/Q _1273_/X _1267_/Y _1473_/Q _1292_/X _1473_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_48_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1005__A _1005_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0844__A _0843_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__B1 _1072_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_37 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1376__A1 _0887_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1376__B2 _1375_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1394__B _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1560__D _1104_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_292 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_67 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0754__A _0728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0920__C _0920_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0929__A _0874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0878__B1 _0870_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_218 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1470__D _1470_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1055__B1 _1537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0814__D _0814_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_170 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1540__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_152 VGND VPWR sky130_fd_sc_hd__fill_2
X_0932_ _0757_/X _1399_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0863_ _0880_/A _0777_/B _0864_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_61_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1563__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_0794_ _1313_/A _0794_/B _0728_/X _1313_/D _0794_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_5_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_1415_ _0885_/A _1415_/B _1415_/C _1415_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__0839__A _0768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_1346_ _0773_/X _1346_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_1277_ _1272_/X _1276_/Y _0707_/B _1241_/X _1277_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1294__B1 _1473_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1389__B _0720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_298 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_36 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1349__A1 _1513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1555__D _1097_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_354 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0828__B1_N _0827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1563__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0931__B _1250_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_144 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0796__C1 _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_166 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1465__D _0806_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_1200_ _1200_/A _1214_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_335 VGND VPWR sky130_fd_sc_hd__decap_8
X_1131_ _1131_/A _1131_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1062_ _1540_/Q _0912_/X _1062_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1276__B1 _0707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1287__A1_N _1272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1002__B _1078_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1291__A3 _1290_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_287 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1028__B1 _0827_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0915_ _0846_/A _0913_/Y _1484_/Q _0914_/Y _0915_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0846_ _0846_/A _0818_/B _0846_/C _0846_/D _0846_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0777_ _0777_/A _0777_/B _0778_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1436__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_346 VGND VPWR sky130_fd_sc_hd__fill_2
X_1329_ _1329_/A _1329_/B _1330_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1586__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_210 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1485__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1019__B1 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_390 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0942__A _0938_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1025__A3 _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0784__A2 _0887_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1459__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_48_A clkbuf_3_7_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1114_ _0920_/C _1150_/B _1114_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_357 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0836__B _0836_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1013__A _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1045_ _0912_/X _0835_/A _0823_/A _0992_/X _1045_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_61_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0852__A _0851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_257 VGND VPWR sky130_fd_sc_hd__fill_2
X_0829_ _0823_/B _0829_/B _0829_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_56_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_357 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_316 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_327 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0762__A _0760_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_22 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1601__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1412__B1 _1409_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1191__A2 _1189_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__A _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_393 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1403__B1 _1350_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1594_ _1218_/X _1217_/A _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1008__A _1536_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_390 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_198 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_179 VGND VPWR sky130_fd_sc_hd__decap_4
X_1028_ _1526_/Q _1018_/X _0827_/B _1021_/X _1028_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_34_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1397__B _1397_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__A2 _0851_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_25 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1563__D _1563_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1173__A2 _1171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0757__A _0756_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0907__D _0907_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_308 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0923__C _1145_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__A2 _0980_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_341 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1473__D _1473_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_249 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1588__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1517__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0978__A2 _0971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_93 VGND VPWR sky130_fd_sc_hd__decap_4
X_1577_ _1168_/X _0916_/A rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_249 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_179 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_116 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_138 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_190 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1201__A _1201_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1558__D _1100_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1146__A2 usb_rst VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_18 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1610__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_282 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1111__A _1560_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_352 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1468__D _1467_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1385__A2 _1397_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1500_ _0954_/X endpoint[3] rst_n _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1431_ _1431_/D data_out[4] _1518_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1362_ _0715_/A _0762_/X _1362_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0896__A1 _1313_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1293_ _1288_/Y _1252_/B _1292_/X _1293_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_55_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1005__B _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_296 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1021__A _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__A1 _0999_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1376__A2 _1400_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1394__C _0869_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_282 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0754__B _0754_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_311 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0770__A _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_78 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_304 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0920__D _1566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1492__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0878__A1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1106__A _0925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0945__A _0754_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_266 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1055__B2 _1016_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0931_ _0874_/C _1250_/A _1300_/A tx_se0 VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_9_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_175 VGND VPWR sky130_fd_sc_hd__decap_4
X_0862_ _0862_/A _0880_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0793_ _0732_/A _1316_/B _1313_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_54_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_311 VGND VPWR sky130_fd_sc_hd__decap_12
X_1414_ _1414_/A _0957_/B _1415_/C VGND VPWR sky130_fd_sc_hd__or2_4
X_1345_ _0772_/C _1339_/X _1330_/A _1344_/Y _1345_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_3_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_366 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1016__A _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1276_ _1421_/Q _1273_/X _0707_/A _1276_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__0855__A _1187_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1294__A1 _1506_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1294__B2 _1292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_274 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1389__C _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1535__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1598__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1349__A2 _0773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1571__D _1144_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_377 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_34 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0765__A _0725_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_11 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_8_0_clk_48_A clkbuf_4_9_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0796__B1 _0794_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0931__C _1300_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1481__D _1291_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_1130_ _0922_/A _1130_/B _1131_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_65_347 VGND VPWR sky130_fd_sc_hd__fill_2
X_1061_ _1016_/X _1060_/X _1539_/Q _1016_/X _1539_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1276__A1 _1421_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_285 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_211 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1028__A1 _1526_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1002__C _1002_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_266 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1028__B2 _1021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_299 VGND VPWR sky130_fd_sc_hd__fill_2
X_0914_ _0910_/X _0914_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0845_ _0851_/D _0846_/D VGND VPWR sky130_fd_sc_hd__inv_8
X_0776_ _0776_/A _0776_/B _0755_/A _0775_/X _0777_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_68_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_174 VGND VPWR sky130_fd_sc_hd__fill_2
X_1328_ _0760_/Y _1326_/X _1315_/A _1327_/X _1328_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_1259_ _1250_/C _0874_/A _1259_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_64_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_406 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1019__A1 _1528_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_14 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1566__D _1125_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_104 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_130 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0950__B1 _0949_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_152 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_141 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1530__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_317 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_266 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_269 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1476__D _1277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0941__B1 _0940_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_369 VGND VPWR sky130_fd_sc_hd__decap_4
X_1113_ _1110_/X _1111_/X _1158_/A _1562_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_65_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40 VGND VPWR sky130_fd_sc_hd__fill_1
X_1044_ _1034_/X _0829_/X _0832_/B _0992_/X _1044_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1013__B _1532_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_394 VGND VPWR sky130_fd_sc_hd__fill_2
X_0828_ _0827_/A _0827_/B _0827_/X _0843_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0759_ _0759_/A _0759_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1553__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14_0_clk_48_A clkbuf_3_7_0_clk_48/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1204__A _1204_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_68 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0762__B _1185_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_12 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1412__A1 _0887_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_29 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1176__B1 _1175_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__B _1492_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_155 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1114__A _0920_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0953__A endpoint[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_309 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1100__B1 _0906_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_372 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1426__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_291 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1403__A1 _1425_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1576__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_1593_ _1593_/D _1593_/Q _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_38_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_1027_ _1020_/X _1037_/A _1018_/A _1525_/Q _0998_/X _1525_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__0863__A _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_372 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0757__B _0757_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1449__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0773__A _0773_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1599__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__A3 _1446_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_70 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1109__A _0919_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_103 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1557__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0877__A2_N _0872_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_331 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0978__A3 _1525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1178__A1_N _0811_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1576_ _1163_/X _1159_/A rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__0858__A _1528_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1312__B1 _1296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_125 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_26 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_342 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1201__B _1604_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_58 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1574__D _1153_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0768__A _0767_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_235 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_261 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1111__B _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_7 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1484__D _1484_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1430_ _1430_/D data_out[3] _1421_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1361_ data_in[0] _1399_/B _1361_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0896__A2 _0794_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1292_ _1247_/D tx_en _0715_/C _1292_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1005__C _1005_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_264 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1302__A _1301_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_128 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1073__A2 _1069_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1376__A3 _1371_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1394__D _1394_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__A1_N _1046_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1559_ _1101_/X _0907_/D rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1212__A _1212_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_106 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0754__C _0862_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1311__B1_N _1310_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1569__D _1135_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_194 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0878__A2 _0865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0945__B _0945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1122__A _1128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1479__D _1283_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0961__A _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0930_ _1194_/B _1250_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0861_ _1358_/A _0861_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0792_ _0776_/B _1316_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_42_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1413_ _0856_/B _1413_/B _1415_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_323 VGND VPWR sky130_fd_sc_hd__decap_12
X_1344_ _0772_/C _1342_/A _1344_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_3_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1572__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_1275_ _1272_/X _1274_/Y _1269_/A _1241_/X _1475_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1501__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1294__A2 _1273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_201 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1389__D _1389_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0871__A _1357_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_256 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1_0_clk_48_A clkbuf_0_clk_48/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_49 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1207__A _1207_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0765__B _0755_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_234 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0781__A data_toggle VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0796__A1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1117__A _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0956__A _1413_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1541__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1060_ _1056_/Y _1059_/Y _1056_/A _1004_/X _1060_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_18_220 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1276__A2 _1273_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_256 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1028__A2 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1002__D _1002_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0913_ _1102_/A _0824_/B _0912_/X _0913_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0844_ _0843_/X _0851_/D VGND VPWR sky130_fd_sc_hd__buf_1
X_0775_ _0774_/X _0775_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0866__A handshake[0] VGND VPWR sky130_fd_sc_hd__diode_2
X_1327_ _0886_/A _1327_/B _1327_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_1258_ _1329_/A _1258_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_1189_ _0718_/X _1189_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_64_392 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_245 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1482__CLK _1609_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_267 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1019__A2 _1016_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_127 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1494__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1582__D _1582_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0950__A1 _1435_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0776__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_337 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_clk_48 clkbuf_3_7_0_clk_48/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_15_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1400__A _1425_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_248 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1492__D _1492_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0941__A1 _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_1112_ _1102_/A _1158_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_348 VGND VPWR sky130_fd_sc_hd__decap_3
X_1043_ _1034_/X _0827_/A _0829_/B _1039_/X _1458_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_0_63 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1013__C _1013_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_381 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_340 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_72 VGND VPWR sky130_fd_sc_hd__decap_4
X_0827_ _0827_/A _0827_/B _0827_/X VGND VPWR sky130_fd_sc_hd__or2_4
Xclkbuf_3_0_0_clk_48 clkbuf_3_1_0_clk_48/A clkbuf_4_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0758_ _0757_/X _0758_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_28_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_315 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_58 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1220__A _1595_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1577__D _1168_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1412__A2 _1407_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1176__A1 _1581_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__C _1313_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1114__B _1150_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_370 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0953__B _0945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1100__B2 _1095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1100__A1 _1557_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1130__A _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1487__D _1487_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1403__A2 _0786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_1592_ _1213_/X _1212_/A _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__1305__A _1305_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_307 VGND VPWR sky130_fd_sc_hd__fill_2
X_1026_ _1020_/X _0834_/B _1018_/A _1524_/Q _0998_/X _1026_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__0863__B _0777_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1520__CLK _1529_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_13 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_115 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_229 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1125__A _1128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1085__B1 _1084_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1543__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1526__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1575_ _1575_/D _1155_/A rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__0858__B _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_207 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1312__B2 tx_j VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0874__A _0874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_310 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VPWR sky130_fd_sc_hd__decap_3
X_1009_ _1536_/Q _0840_/X _1008_/Y _0841_/Y _1009_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_22_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1590__D _1590_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1566__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_118 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_310 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clk_48 clkbuf_4_3_0_clk_48/A _1518_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1111__C _0919_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1360_ transaction_active _1359_/X _1329_/B _1360_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA_clkbuf_2_3_0_clk_48_A clkbuf_2_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_280 VGND VPWR sky130_fd_sc_hd__fill_2
X_1291_ _1288_/Y _1267_/Y _1290_/X _1285_/Y _1241_/X _1291_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_36_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_251 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1005__D _1004_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_295 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_232 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1058__B1 _1537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1439__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0869__A _0869_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1558_ _1100_/X _0906_/A rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1489_ _0765_/X _0724_/A rst_n _1577_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1589__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1212__B _1214_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0754__D _0754_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1049__B1 _1532_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1585__D _1179_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1221__B1 _1220_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0779__A _0779_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_402 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1122__B _1122_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_224 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_0860_ _0732_/A _0856_/X _1413_/B _0879_/B VGND VPWR sky130_fd_sc_hd__o21a_4
X_0791_ _0791_/A _0794_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1495__D _1495_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1412_ _0887_/A _1407_/X _1409_/Y _1411_/X _1412_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_68_335 VGND VPWR sky130_fd_sc_hd__decap_6
X_1343_ _0772_/A _0772_/B _1330_/X _1342_/Y _1510_/D VGND VPWR sky130_fd_sc_hd__a211o_4
X_1274_ _1420_/Q _1273_/X _0707_/B _1274_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1279__B1 _0707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1313__A _1313_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1294__A3 _1267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_279 VGND VPWR sky130_fd_sc_hd__fill_2
X_0989_ _0901_/A _0970_/X _0744_/B data_out[5] _0961_/X _0989_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_59_324 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0765__C _0764_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_46 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1604__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0796__A2 _0790_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_158 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1117__B _0920_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0972__A _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1054__A1_N _1008_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0912_ _0818_/B _0912_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0843_ _0843_/A _0843_/B _0843_/C _0842_/Y _0843_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0774_ _1513_/Q _0773_/X _0774_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1308__A _1301_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_121 VGND VPWR sky130_fd_sc_hd__decap_3
X_1326_ _0869_/A _0725_/B _1327_/B _1326_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_68_187 VGND VPWR sky130_fd_sc_hd__fill_2
X_1257_ _1241_/X _1255_/X _1256_/X _1257_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_17_39 VGND VPWR sky130_fd_sc_hd__fill_2
X_1188_ _1470_/Q _1185_/B _1186_/Y _1187_/X _1470_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_117 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1188__C1 _1187_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0831__A1_N _0829_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0950__A2 _0942_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0776__B _0776_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_235 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0792__A _0776_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1400__B _1400_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_82 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1128__A _1128_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0941__A2 _0945_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_327 VGND VPWR sky130_fd_sc_hd__decap_4
X_1111_ _1560_/Q _0919_/B _0919_/C _1150_/B _1111_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_48_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_157 VGND VPWR sky130_fd_sc_hd__decap_4
X_1042_ _1034_/X _0837_/X _0825_/B _1039_/X _1042_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_46_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_95 VGND VPWR sky130_fd_sc_hd__fill_2
X_0826_ _0994_/A _0826_/B _0827_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_0757_ _0756_/Y _0757_/B _0757_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_29_349 VGND VPWR sky130_fd_sc_hd__fill_2
X_1309_ _1309_/A _1309_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_44_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_363 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1220__B _1222_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_238 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1593__D _1593_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1176__A2 _1171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0787__A _1381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1100__A2 _1090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1130__B _1130_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_242 VGND VPWR sky130_fd_sc_hd__fill_2
X_1591_ _1591_/D _1591_/Q _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_7_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_80 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1472__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_102 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1305__B _1305_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_127 VGND VPWR sky130_fd_sc_hd__fill_2
X_1025_ _1020_/X _0836_/B _1018_/A _1523_/Q _1021_/X _1523_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_34_352 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1321__A _0780_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1328__A2_N _1326_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0809_ _0808_/X _1102_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_330 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1588__D _0768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_clk_48_A clkbuf_3_5_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1251__D1 _1250_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1495__CLK _1577_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1406__A _1406_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1125__B _1125_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1141__A _0918_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_330 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1085__A1 _1002_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1498__D _1498_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0980__A _0970_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_355 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_399 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1566__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VPWR sky130_fd_sc_hd__fill_2
X_1574_ _1153_/X _1154_/A rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1316__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0874__B _0874_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1051__A _1014_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_149 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VPWR sky130_fd_sc_hd__decap_3
X_1008_ _1536_/Q _1008_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_41_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0890__A _0777_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_366 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1226__A _1598_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_274 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_344 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1111__D _1150_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_399 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1136__A _0918_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_270 VGND VPWR sky130_fd_sc_hd__fill_2
X_1290_ _1289_/Y _1247_/D _1290_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_0_292 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1510__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1058__B2 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_174 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0869__B _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1557_ _1557_/D _1557_/Q rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1046__A _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0741__B1 usb_address[3] VGND VPWR sky130_fd_sc_hd__diode_2
X_1488_ _1488_/D _1358_/A rst_n _1514_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_39_252 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0885__A _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_296 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1049__B2 _1036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1221__A1 _1217_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1533__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__A _0715_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_189 VGND VPWR sky130_fd_sc_hd__fill_2
X_0790_ _0887_/B _0786_/Y _0786_/Y _0789_/X _0790_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1411_ _0769_/Y _0725_/B _1406_/A _1410_/X _1411_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_303 VGND VPWR sky130_fd_sc_hd__decap_6
X_1342_ _1342_/A _1342_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_3_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_86 VGND VPWR sky130_fd_sc_hd__fill_2
X_1273_ _1269_/B _1273_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1279__B2 _1240_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1313__B _0879_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_244 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_266 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1299__A1_N _1201_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_225 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1581__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1510__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_0988_ _0901_/A _0970_/X _1447_/Q data_out[4] _0961_/X _1431_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1237__A1_N _1236_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1556__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_1609_ _1609_/D _0873_/A rst_n _1609_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_358 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1596__D _1596_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_144 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_84 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1117__C _0925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_306 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1414__A _1414_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1429__CLK _1421_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0911_ _0818_/X _0901_/Y _1484_/Q _0910_/X _1484_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1579__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0842_ _0837_/X _0841_/Y _0837_/X _0841_/Y _0842_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
X_0773_ _0773_/A _0773_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_52_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0944__B1 _0943_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1308__B _1307_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_133 VGND VPWR sky130_fd_sc_hd__fill_2
X_1325_ _0867_/B _1321_/Y _1324_/X _1325_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_56_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1324__A _1324_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1256_ _1245_/X _1252_/B _1250_/A _1256_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_1187_ _1187_/A _1187_/B _1187_/C _1187_/X VGND VPWR sky130_fd_sc_hd__or3_4
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1188__B1 _1186_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1234__A _1234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0776__C _0755_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_306 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1360__B1 _1329_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_394 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1409__A _1409_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1179__B1 _0814_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1128__B _1128_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1351__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1110_ _1109_/Y _1107_/Y _1110_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1144__A _1158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1103__B1 _1560_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VPWR sky130_fd_sc_hd__fill_2
X_1041_ _1034_/X _0835_/B _0836_/B _1039_/X _1456_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_46_350 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_353 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1319__A _1319_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0825_ _0821_/Y _0825_/B _0827_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_0756_ data_in_valid _0756_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_4_7_0_clk_48_A clkbuf_4_7_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_1308_ _1301_/X _1307_/X _1612_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0893__A _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1239_ _1214_/B _1238_/X _1604_/Q _1205_/X _1239_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_52_331 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_26 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1053__A1_N _1014_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_342 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_397 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1139__A _0925_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1590_ _1590_/D _1207_/A _0928_/X _1466_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_15_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1305__C _0712_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_136 VGND VPWR sky130_fd_sc_hd__fill_2
X_1024_ _1020_/X _0825_/B _1018_/X _1522_/Q _1021_/X _1024_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_19_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_331 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1321__B _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_0808_ _0808_/A _0808_/B _0808_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_0739_ usb_address[2] _0738_/Y _0739_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_29_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_194 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1251__C1 _1248_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0798__A _0798_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1406__B _1362_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_82 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13_0_clk_48_A clkbuf_3_6_0_clk_48/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1085__A2 _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_378 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_64 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1547__SET_B _0927_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1573_ _1573_/D _1573_/Q rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1316__B _1316_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0874__C _0874_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1051__B _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1007_ _0791_/A _0996_/X _1006_/X _1530_/D VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_22_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_28 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1226__B _1222_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_286 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1242__A _0874_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1599__D _1229_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_40 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1462__CLK _1466_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_83 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1312__A2_N _1296_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_242 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1152__A _1154_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_256 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1327__A _0886_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1556_ _1098_/X _1556_/Q rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__0741__B2 _0740_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1487_ _1487_/D _0777_/A rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__0885__B _0884_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1062__A _1540_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_245 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1485__CLK _1472_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_304 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_308 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1221__A2 _1216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1405__A1_N _1401_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1593__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__B _1185_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_142 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1147__A _1147_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1410_ _1350_/X _1410_/B _1410_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_1341_ _1340_/X _1342_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1272_ _1272_/A _1272_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_201 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1313__C _1315_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_19 VGND VPWR sky130_fd_sc_hd__fill_1
X_0987_ _0979_/X _0980_/X _1446_/Q data_out[3] _0981_/X _1430_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1057__A _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1608_ _1257_/Y _0874_/A rst_n _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1603__SET_B _0928_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1539_ _1539_/D _1539_/Q _0927_/X _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_47_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_256 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_63 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1500__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1414__B _0957_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_0910_ _0909_/X _0910_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0841_ _0840_/X _0841_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0772_ _0772_/A _0772_/B _0772_/C _1512_/Q _0773_/A VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0944__A1 _0755_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_112 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_1324_ _1324_/A _1323_/X _1324_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_156 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_318 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1324__B _1323_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1255_ _1252_/A _1196_/A _1254_/X _1255_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1121__A1 _0920_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1186_ _1186_/A _1186_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1340__A _1339_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1523__CLK _1443_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1188__A1 _1470_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1234__B _1200_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0776__D _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1360__A1 transaction_active VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1250__A _1250_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1283__A1_N _1272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1409__B _1409_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1179__B2 _1092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1179__A1 _0811_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_0_0_clk_48_A clkbuf_0_clk_48/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1351__A1 _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1144__B _1144_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22 VGND VPWR sky130_fd_sc_hd__fill_1
X_1040_ _1034_/X _0830_/X _0834_/B _1039_/X _1040_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1103__B2 usb_rst VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_373 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1160__A _1160_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1546__CLK _1454_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_292 VGND VPWR sky130_fd_sc_hd__fill_2
X_0824_ _1187_/C _0824_/B _0846_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1319__B _1318_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0755_ _0755_/A _0755_/B _1329_/B _0755_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__1335__A _1509_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_137 VGND VPWR sky130_fd_sc_hd__fill_2
X_1307_ _1612_/Q _1306_/B _1612_/Q _1306_/B _1307_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_159 VGND VPWR sky130_fd_sc_hd__fill_2
X_1238_ _1603_/Q _1204_/Y _1236_/Y _1204_/A _1238_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_1169_ _0916_/C _1165_/X _1158_/A _1578_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1070__A _0999_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_207 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_49 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1030__B1 _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1419__CLK _1514_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1245__A _0874_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1569__CLK _1575_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1097__B1 _1555_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_332 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_50 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_200 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1139__B _1138_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1155__A _1155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0994__A _0994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_159 VGND VPWR sky130_fd_sc_hd__fill_2
X_1023_ _1020_/X _0829_/B _1018_/X _1521_/Q _1021_/X _1521_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1088__B1 _1086_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_19 VGND VPWR sky130_fd_sc_hd__decap_4
X_0807_ _0797_/Y _0803_/X _0806_/Y _0808_/B VGND VPWR sky130_fd_sc_hd__o21a_4
X_0738_ _1445_/Q _0738_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1065__A _1001_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_49 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1079__B1 _1078_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_357 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1251__B1 _1247_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__A1_N _0747_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_107 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_clk_48 clkbuf_2_1_0_clk_48/A clkbuf_3_1_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_32 VGND VPWR sky130_fd_sc_hd__decap_4
X_1572_ _1572_/D _1145_/A rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_3_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1575__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1504__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_170 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_1006_ _0998_/X _1006_/B _1006_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_22_346 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_390 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1233__B1 _1232_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__A _1358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1607__CLK _1589_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1152__B _1150_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_268 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1215__B1 _1214_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1327__B _1327_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1555_ _1097_/X _1555_/Q rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1486_ _0915_/X _0901_/B rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1062__B _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1206__B1 _1589_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_198 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1497__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__C _0724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_61 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1147__B _1149_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1340_ _1339_/X _1340_/B _1340_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_3_33 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_66 VGND VPWR sky130_fd_sc_hd__fill_1
X_1271_ _1267_/Y _1269_/X _1270_/X _1201_/A _1240_/X _1271_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1133__C1 _1132_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1313__D _1313_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_238 VGND VPWR sky130_fd_sc_hd__fill_2
X_0986_ _0979_/X _0980_/X _1445_/Q data_out[2] _0981_/X _0986_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_1607_ _1607_/D _0874_/B rst_n _1589_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xclkbuf_3_3_0_clk_48 clkbuf_3_3_0_clk_48/A clkbuf_4_7_0_clk_48/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1538_ _1538_/D _1056_/A _0927_/X _1529_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1469_ _0766_/A _0766_/B _1467_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1452__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_28 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_202 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_2_0_clk_48_A clkbuf_2_3_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_113 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_102 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1248__A _1250_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1607__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_0840_ _0838_/Y _0768_/X _1461_/Q _1187_/B _0840_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_0771_ _0771_/A _0771_/B _1509_/Q _0772_/B VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1158__A _1158_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1475__CLK _1611_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_161 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0944__A2 _0941_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0997__A _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1323_ _0861_/Y _0778_/B _0795_/X _1322_/X _1323_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_1254_ _0874_/A _1252_/A _0874_/C _1254_/D _1254_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_49_382 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_330 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1121__A2 _1117_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1185_ _1470_/Q _1185_/B _1186_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_64_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1340__B _1340_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_249 VGND VPWR sky130_fd_sc_hd__fill_1
X_0969_ _1187_/A _0969_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1188__A2 _1185_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1345__C1 _1344_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1360__A2 _1359_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1250__B _1245_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_219 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_400 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1498__CLK _1518_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1409__C _1408_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1179__A2 _1090_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1351__A2 _0789_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_308 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1144__C _1143_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67 VGND VPWR sky130_fd_sc_hd__fill_1
X_0823_ _0823_/A _0823_/B _0824_/B VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__1529__RESET_B rst_n VGND VPWR sky130_fd_sc_hd__diode_2
X_0754_ _0728_/X _0754_/B _0862_/A _0754_/D _1329_/B VGND VPWR sky130_fd_sc_hd__nor4_4
X_1306_ _1304_/Y _1306_/B _1301_/X _1306_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_56_116 VGND VPWR sky130_fd_sc_hd__decap_4
X_1237_ _1236_/Y _1208_/X _1234_/A _1208_/X _1237_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_1168_ _0916_/C _1166_/Y _1147_/A _1167_/X _1168_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_52_311 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1070__B _1064_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1501__D _0946_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1099_ _1556_/Q _1094_/X _1557_/Q _1095_/X _1557_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_20_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1030__B2 _0853_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1030__A1 _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_105 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_341 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1097__A1 _1554_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1097__B2 _1095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_363 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_374 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_73 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_clk_48 clkbuf_4_7_0_clk_48/A _1472_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1155__B _1155_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_81 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1513__CLK _1467_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0994__B _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1022_ _1020_/X _0832_/B _1018_/X _1520_/Q _1021_/X _1022_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1088__B2 _1004_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1088__A1 _1086_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_300 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1171__A _1092_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0806_ _0806_/A _0805_/X _0806_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0737_ _0856_/B _1313_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1346__A _0773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1065__B _1064_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_17 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1079__A1 _1002_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_369 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1251__A1 _1252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_226 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1536__CLK _1583_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_366 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_83 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1571_ _1144_/Y _0918_/A rst_n _1575_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__1166__A _1165_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_119 VGND VPWR sky130_fd_sc_hd__decap_4
X_1005_ _1005_/A _1001_/X _1005_/C _1004_/X _1006_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_19_193 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_358 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1233__A1 _1600_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1559__CLK _1567_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__B _0892_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1076__A _1002_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1049__A2_N _1036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_314 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_144 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0983__B1 _1442_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__B1 usb_address[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_299 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1215__A1 _1212_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0974__B1 _1436_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1554_ _1554_/D _1554_/Q rst_n _1567_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_3_4_0_clk_48_A clkbuf_3_5_0_clk_48/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1485_ _0847_/X _1485_/Q rst_n _1472_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
.ends


* NGSPICE file created from usb_cdc_core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 D Q RESET_B CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 D Q SET_B CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 Y VGND VPWR
.ends

.subckt usb_cdc_core clk_i enable_i inport_accept_o inport_data_i[0] inport_data_i[1]
+ inport_data_i[2] inport_data_i[3] inport_data_i[4] inport_data_i[5] inport_data_i[6]
+ inport_data_i[7] inport_valid_i outport_accept_i outport_data_o[0] outport_data_o[1]
+ outport_data_o[2] outport_data_o[3] outport_data_o[4] outport_data_o[5] outport_data_o[6]
+ outport_data_o[7] outport_valid_o rst_i utmi_data_in_i[0] utmi_data_in_i[1] utmi_data_in_i[2]
+ utmi_data_in_i[3] utmi_data_in_i[4] utmi_data_in_i[5] utmi_data_in_i[6] utmi_data_in_i[7]
+ utmi_data_out_o[0] utmi_data_out_o[1] utmi_data_out_o[2] utmi_data_out_o[3] utmi_data_out_o[4]
+ utmi_data_out_o[5] utmi_data_out_o[6] utmi_data_out_o[7] utmi_dmpulldown_o utmi_dppulldown_o
+ utmi_linestate_i[0] utmi_linestate_i[1] utmi_op_mode_o[0] utmi_op_mode_o[1] utmi_rxactive_i
+ utmi_rxerror_i utmi_rxvalid_i utmi_termselect_o utmi_txready_i utmi_txvalid_o utmi_xcvrselect_o[0]
+ utmi_xcvrselect_o[1] VPWR VGND
XANTENNA__4357__D _3362_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_222 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_19 VGND VPWR sky130_fd_sc_hd__fill_1
X_3155_ _3219_/A _3014_/Y _3088_/Y _3158_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_27_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_545 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3086_ _3015_/X _3360_/A _3071_/A _3105_/D _3086_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2455__A _2456_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2651__B1 _4522_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2977__A2_N _2976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_689 VGND VPWR sky130_fd_sc_hd__fill_2
X_3988_ _3987_/Y _3979_/X _3929_/Y _3981_/X _3988_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2902__B _3491_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2939_ _2938_/X _2940_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_486 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_328 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3286__A _3243_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4490__RESET_B _2307_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2190__A _2188_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4609_ _4609_/D _4236_/A _2164_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_422 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3903__B1 _3902_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_66 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_444 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_433 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_199 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_520 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3131__A1 _3085_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_501 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_383 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_545 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2890__B1 _2996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_214 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2365__A _2362_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4092__C1 _4091_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_475 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4578__RESET_B _2201_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_667 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3908__B _3904_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4507__RESET_B _2286_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_148 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3198__A1 _3019_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2812__B _2799_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3196__A _3031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2531__C _2528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_310 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_230 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3643__B _3640_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3370__A1 _3369_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_626 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3362__C _3362_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_582 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_203 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2275__A _2277_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2881__B1 _2871_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_397 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_589 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2706__C _2562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4193__C _4192_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_91 VGND VPWR sky130_fd_sc_hd__fill_2
X_3911_ _3005_/Y _2560_/X _3911_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3842_ _4530_/Q _3830_/X _3842_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_615 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3818__B _3804_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_497 VGND VPWR sky130_fd_sc_hd__fill_2
X_3773_ _3769_/X _3772_/X _3720_/A _3773_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_2724_ _2724_/A _2544_/X _2724_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_569 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_2655_ _2680_/A _2654_/X _2655_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_192 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3834__A _4519_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3553__B _3541_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4400__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_604 VGND VPWR sky130_fd_sc_hd__fill_2
X_4325_ _3323_/Y _2909_/A _2504_/X _4325_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2586_ _2560_/X _3417_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_637 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_615 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_339 VGND VPWR sky130_fd_sc_hd__fill_2
X_4256_ _4232_/Y _4263_/B _4258_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_95_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_361 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_4187_ _4137_/B _4146_/B _4187_/C _4187_/D _4187_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_3207_ _3207_/A _3199_/Y _3207_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_715 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4550__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3664__A2 _3430_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3138_ _3227_/D _3095_/X _3138_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_27_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_353 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_707 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_68 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_589 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4074__C1 _4073_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2185__A _2183_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3069_ _3046_/X _3038_/Y _3011_/X _3010_/X _3069_/X VGND VPWR sky130_fd_sc_hd__or4_4
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2913__A _3319_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_615 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_475 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4600__RESET_B _2176_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4550__D _3907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3463__B _3463_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_346 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4278__C _4278_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_350 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4301__B1 _4300_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_203 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2807__B _2666_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_556 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_258 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_526 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2526__C _2526_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_559 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_537 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2823__A _2796_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_250 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3919__A _4318_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4080__A2 _4056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3638__B _3625_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4341__RESET_B _2485_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_497 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4460__D _4522_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4423__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_528 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3654__A _3554_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2440_ _2443_/A _2440_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_108_591 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3343__A1 _3330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3894__A2 _3883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_615 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4188__C _4188_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2371_ _2367_/X _2371_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_648 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4573__CLK _4574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4110_ _3915_/Y _4562_/Q _3915_/Y _4562_/Q _4110_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_618 VGND VPWR sky130_fd_sc_hd__fill_2
X_4041_ _4041_/A _4039_/B _4041_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_94_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_180 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_206 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4429__RESET_B _2379_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_280 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2733__A _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3548__B _3546_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_592 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_581 VGND VPWR sky130_fd_sc_hd__fill_2
X_3825_ _3824_/X _3904_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4370__D _3662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_311 VGND VPWR sky130_fd_sc_hd__fill_2
X_3756_ _2658_/Y _2659_/X _4525_/Q _2650_/Y _3759_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2947__A1_N _4428_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2707_ _2707_/A _2706_/X _2707_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3687_ _3687_/A _3687_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3564__A _3506_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2638_ _3704_/A _2638_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3885__A2 _3883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_250 VGND VPWR sky130_fd_sc_hd__fill_2
X_2569_ _2568_/B _2562_/X _2566_/X _2705_/B _2569_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_59_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_4308_ _4247_/A _2707_/A _4307_/Y _4308_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_101_266 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_629 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_169 VGND VPWR sky130_fd_sc_hd__fill_2
X_4239_ _4234_/Y _4368_/Q _4249_/A _4238_/X _4239_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_101_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2908__A _2886_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_320 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2845__B1 _2844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_534 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4545__D _3896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_312 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4047__C1 _4046_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_548 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3739__A _3671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2643__A _4520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_378 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_48 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3458__B _3458_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_261 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4446__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_311 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_449 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3177__C _3097_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3474__A _3483_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4596__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_622 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_110 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3193__B _3186_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_520 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3876__A2 _3869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_594 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2818__A _2818_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3089__B1 _3055_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_512 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_448 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2537__B _3818_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_556 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4455__D _2671_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_375 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4593__RESET_B _2184_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4522__RESET_B _2269_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3649__A _3581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_209 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3800__A2 _3785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4109__B1_N _4108_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2553__A _4620_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_66 VGND VPWR sky130_fd_sc_hd__decap_3
X_3610_ _4392_/Q _3610_/B _3610_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3365__B1_N _3369_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4590_ _4590_/D _4185_/A _2187_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3541_ _3513_/A _3541_/B _3542_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3384__A _3397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_347 VGND VPWR sky130_fd_sc_hd__decap_12
X_3472_ _3486_/B _3479_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3316__A1 _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4199__B _4199_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2423_ _2419_/A _2423_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3316__B2 _3248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_412 VGND VPWR sky130_fd_sc_hd__decap_6
X_2354_ _2358_/A _2354_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3831__B _3830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_618 VGND VPWR sky130_fd_sc_hd__fill_2
X_2285_ _2283_/A _2285_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2728__A _4500_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4319__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_459 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2827__B1 _2783_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_320 VGND VPWR sky130_fd_sc_hd__fill_2
X_4024_ _4564_/Q _4024_/B _4024_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4365__D _3401_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4292__A2 _4284_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_353 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_559 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3559__A _3559_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_676 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4469__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_209 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4044__A2 _4037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_36 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_25 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2463__A _2460_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3808_ _3808_/A _3805_/X _3808_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3004__B1 _2996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_697 VGND VPWR sky130_fd_sc_hd__decap_4
X_3739_ _3671_/X _3739_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3294__A _3243_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2910__B _2910_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_38 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_614 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2638__A _3704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_407 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_97 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3469__A _3498_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_367 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4035__A2 _4034_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2373__A _2367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_581 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3794__B2 _3792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3794__A1 _2684_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3188__B _3220_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_703 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_275 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_130 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4095__B1_N _4094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_485 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3651__B _3646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_82 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2548__A _2548_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4611__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_301 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_676 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_654 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3379__A _3317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2283__A _2283_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2972_ _2972_/A _2972_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_91_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2730__B _4504_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4573_ _4092_/X _3947_/A _2207_/X _4574_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__3545__C _3545_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_634 VGND VPWR sky130_fd_sc_hd__decap_6
X_3524_ _2863_/B _3513_/B _3524_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_103_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_3455_ _3455_/A _3434_/B _3458_/B VGND VPWR sky130_fd_sc_hd__nor2_4
X_2406_ _2408_/A _2406_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3842__A _4530_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_562 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3561__B _3582_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_253 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_231 VGND VPWR sky130_fd_sc_hd__fill_2
X_3386_ _3385_/X _3386_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_350 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_2337_ _2337_/A _2337_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2458__A _2456_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_106 VGND VPWR sky130_fd_sc_hd__fill_2
X_2268_ _2272_/A _2268_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4444__RESET_B _2362_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_407 VGND VPWR sky130_fd_sc_hd__decap_12
X_4007_ _4007_/A _4007_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_53_632 VGND VPWR sky130_fd_sc_hd__fill_1
X_2199_ _2199_/A _2199_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_35 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3289__A _3289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2905__B _4418_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_186 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2193__A _2188_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3776__B2 _3771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2921__A _2920_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3736__B _3734_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2640__B _3707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_166 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3174__D _3173_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3471__B _3478_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_562 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3700__B2 _3699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_466 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2368__A _2367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_245 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4286__C _4285_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3190__C _3190_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_204 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_654 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3199__A _3087_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_495 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_315 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_326 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3927__A _4319_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_573 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_83 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2831__A _2829_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_595 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3646__B _3528_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2990__A2 _2986_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2550__B _2549_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_304 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2742__A2 _2741_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3662__A _3662_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_271 VGND VPWR sky130_fd_sc_hd__fill_2
X_3240_ _3240_/A _3268_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2278__A _2277_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3381__B _3376_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_415 VGND VPWR sky130_fd_sc_hd__fill_2
X_3171_ _3171_/A _3171_/B _3130_/X _3171_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_86_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2709__C _4502_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_565 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_481 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2725__B _4488_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_643 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_315 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3837__A _3837_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2955_ _2954_/Y _4418_/Q _2954_/Y _4418_/Q _2955_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__4507__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2886_ _4375_/Q _2884_/Y _2896_/A _2886_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__2741__A _2718_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_381 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3556__B _3556_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4556_ _4556_/D _4556_/Q _2228_/X _4619_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4183__A1 _4182_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4183__B2 _4180_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3507_ _3504_/A _3505_/Y _3507_/C _3507_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_116_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3930__A1 _2604_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_615 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3572__A _3508_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_315 VGND VPWR sky130_fd_sc_hd__fill_2
X_4487_ _3787_/X _4487_/Q _2311_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3930__B2 _3929_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_13 VGND VPWR sky130_fd_sc_hd__fill_2
X_3438_ _3424_/X _3434_/Y _3437_/X _4426_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_58_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_3369_ _3369_/A _3369_/B _3369_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2188__A _2166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3694__B1 _3687_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_418 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_407 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2916__A _2915_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_462 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_602 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4553__D _4553_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_359 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3747__A _3746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_178 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3466__B _3462_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_475 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3482__A _3513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4366__RESET_B _2455_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_478 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_543 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_296 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_237 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_72 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2826__A _2825_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_568 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_643 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3988__A1 _3987_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3988__B2 _3981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4463__D _4525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4021__A2_N _4020_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_613 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_270 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_646 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_657 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3657__A _2763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3079__D _4355_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_668 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VPWR sky130_fd_sc_hd__decap_3
X_2740_ _2713_/X _2731_/X _2730_/X _2740_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__2561__A _2560_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2671_ _2671_/A _2669_/X _2670_/X _2671_/D _4508_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_4410_ _4410_/D _4410_/Q _2402_/X _4410_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_412 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_646 VGND VPWR sky130_fd_sc_hd__decap_4
X_4341_ _3317_/Y _3314_/A _2485_/X _4430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3392__A _3392_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4272_ _4234_/Y _4253_/A _4272_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_113_489 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_106 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_329 VGND VPWR sky130_fd_sc_hd__decap_6
X_3223_ _3085_/A _3223_/B _3224_/D VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_79_381 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4473__SET_B _2327_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_554 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_3154_ _3059_/Y _3080_/Y _3085_/B _3154_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_94_373 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2736__A _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_289 VGND VPWR sky130_fd_sc_hd__fill_2
X_3085_ _3085_/A _3085_/B _3208_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_27_418 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_248 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_12_0_clk_i clkbuf_3_6_0_clk_i/X clkbuf_5_25_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__4373__D _3422_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_462 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_590 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2651__B2 _2650_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2651__A1 _2649_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_657 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3567__A _3510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_307 VGND VPWR sky130_fd_sc_hd__decap_3
X_3987_ _3987_/A _3987_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2938_ _3302_/A _2979_/A _2938_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2471__A _2472_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2902__C _3494_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3286__B _2973_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_228 VGND VPWR sky130_fd_sc_hd__fill_1
X_2869_ _4379_/Q _2869_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4608_ _4608_/D _4608_/Q _2165_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_2_506 VGND VPWR sky130_fd_sc_hd__decap_12
X_4539_ _3882_/X _4539_/Q _2248_/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3903__A1 _3884_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_78 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4548__D _3903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3131__A2 _3066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_684 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2646__A _2645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2890__A1 _2852_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3828__A2_N _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4092__B1 _4033_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_657 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_167 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3477__A _3483_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2381__A _2381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_127 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3198__A2 _3107_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_690 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3196__B _3360_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4547__RESET_B _2239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2531__D _2531_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_272 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3370__A2 _3369_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_242 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4458__D _4520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3658__B1 _3585_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_510 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_594 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_384 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2881__A1 _2878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_524 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2556__A _4489_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_708 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4352__CLK _4325_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_376 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2706__D _2587_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_473 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_281 VGND VPWR sky130_fd_sc_hd__fill_2
X_3910_ _4317_/Q _2585_/A _3910_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_17_484 VGND VPWR sky130_fd_sc_hd__decap_4
X_3841_ _3883_/A _3841_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3772_ _3695_/B _3771_/X _3695_/B _3771_/X _3772_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_3 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2291__A _2288_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3387__A _3386_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_650 VGND VPWR sky130_fd_sc_hd__fill_2
X_2723_ _2707_/X _2722_/Y _2602_/X _2723_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_9_672 VGND VPWR sky130_fd_sc_hd__fill_2
X_2654_ _2642_/X _2654_/B _2654_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3834__B _3830_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2585_ _2585_/A _3960_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_432 VGND VPWR sky130_fd_sc_hd__decap_12
X_4324_ _4324_/D _4324_/Q _2505_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4011__A utmi_data_out_o[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_415 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_487 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4368__D _3412_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_649 VGND VPWR sky130_fd_sc_hd__fill_1
X_4255_ _4265_/A _4252_/X _4254_/Y _4255_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_101_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_4186_ _4164_/Y _4186_/B _4186_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3206_ _3350_/C _3359_/B _3031_/X _3114_/X _3206_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_55_513 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2466__A _2460_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3137_ _3137_/A _3207_/A _3136_/X _3137_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_55_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_237 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_719 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4074__B1 _4050_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3068_ _3067_/X _3068_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_82_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3821__B1 _3820_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_410 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2913__B _2913_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_605 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3297__A _3297_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_627 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_498 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_504 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_108 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_137 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_44 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_15 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3888__B1 _3887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3463__C _3462_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4278__D _4278_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3760__A _3708_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4375__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4301__A1 _4292_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2376__A _2379_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_492 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2807__C _2805_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_708 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2823__B _2818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3919__B _2585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3000__A _4231_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3935__A _4320_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_660 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4381__RESET_B _2437_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_642 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_631 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_682 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_570 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3654__B _3646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_581 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3343__A2 _3340_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_413 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_627 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4188__D _4188_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2370_ _2367_/X _2370_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3670__A _3705_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_159 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_391 VGND VPWR sky130_fd_sc_hd__fill_2
X_4040_ _4562_/Q _4037_/X _4033_/X _4039_/Y _4562_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_83_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2286__A _2283_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_708 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_22_0_clk_i_A clkbuf_5_22_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_229 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4469__RESET_B _2332_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2733__B _2727_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_3824_ _3824_/A utmi_rxvalid_i _3824_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3548__C _3547_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_446 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_3755_ _3726_/X _3713_/B _3719_/X _3754_/X _4481_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_118_356 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3845__A _4531_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3686_ _2646_/Y _3685_/X _2676_/X _3687_/A VGND VPWR sky130_fd_sc_hd__o21a_4
X_2706_ _2706_/A _2910_/B _2562_/X _2587_/Y _2706_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_106_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3564__B _3582_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2637_ _4447_/Q _3704_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4398__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_540 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_262 VGND VPWR sky130_fd_sc_hd__fill_2
X_2568_ _2580_/A _2568_/B _2705_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_2499_ _2497_/A _2499_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3580__A _3522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_284 VGND VPWR sky130_fd_sc_hd__fill_2
X_4307_ _2706_/X _4307_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_101_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_619 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_159 VGND VPWR sky130_fd_sc_hd__decap_3
X_4238_ _4236_/Y _4260_/A _4237_/Y _4270_/A _4238_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_289 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_660 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2908__B _2906_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4295__B1 _4247_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2196__A _2199_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2845__A1 _4323_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4169_ _4188_/C _4167_/B _4169_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_546 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_708 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4047__B1 _4033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2924__A _4331_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_527 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_582 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_571 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4561__D _4561_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_273 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3458__C _3457_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_457 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_367 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3474__B _3471_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_133 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3193__C _3193_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_435 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_554 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3490__A _3504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3089__A1 _3043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_438 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2818__B _2799_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_524 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2537__C _4501_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_674 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2834__A inport_data_i[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_335 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_387 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3649__B _3649_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4471__D _4471_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3800__A3 _4496_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_34 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2553__B utmi_txready_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_593 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_295 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_93 VGND VPWR sky130_fd_sc_hd__decap_6
X_3540_ _4405_/Q _3543_/B _3542_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4540__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3665__A _4469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2772__B1 _4612_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3384__B _3380_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_450 VGND VPWR sky130_fd_sc_hd__decap_8
X_3471_ _4418_/Q _3478_/B _3471_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_359 VGND VPWR sky130_fd_sc_hd__decap_6
X_2422_ _2419_/A _2422_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3316__A2 _3314_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_221 VGND VPWR sky130_fd_sc_hd__fill_2
X_2353_ _2339_/A _2358_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_565 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_479 VGND VPWR sky130_fd_sc_hd__decap_4
X_2284_ _2283_/A _2284_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4023_ _3969_/Y utmi_data_out_o[7] _3969_/Y _3976_/X _4024_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__2827__A1 _4467_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_516 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_324 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2744__A _4468_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3559__B _3566_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_688 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4381__D _3633_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_582 VGND VPWR sky130_fd_sc_hd__fill_2
X_3807_ _2643_/Y _3803_/X _3806_/X _3807_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3004__A1 _2999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3575__A _3581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_276 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_315 VGND VPWR sky130_fd_sc_hd__fill_2
X_3738_ _3726_/X _3675_/B _3719_/X _3737_/Y _3738_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3294__B _2946_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3669_ _3683_/A _4474_/Q _3669_/C _3668_/X _3669_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_106_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_329 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_318 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3712__C1 _3711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2919__A _2918_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_107 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4556__D _4556_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_10 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_630 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_460 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4413__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2654__A _2642_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_549 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3779__C1 _3778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3469__B _3528_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_20 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_699 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_571 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3794__A2 _3782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3188__C _3188_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4563__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_203 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3485__A _2900_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2754__B1 _2753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3703__C1 _3702_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2829__A _2829_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_392 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_351 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2809__A1 _4514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4466__D _2783_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_354 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_611 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_313 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2564__A _2705_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_666 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3379__B _3379_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_368 VGND VPWR sky130_fd_sc_hd__decap_4
X_2971_ _2953_/Y _2964_/X _2967_/Y _2970_/Y _2971_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_61_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_92 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3395__A _3386_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_585 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2730__C _2729_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4572_ _4086_/X _3939_/A _2208_/X _4574_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_116_646 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_112 VGND VPWR sky130_fd_sc_hd__fill_2
X_3523_ _3514_/A _3521_/Y _3523_/C _3523_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_6_280 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_3454_ _3424_/X _3451_/Y _3453_/X _3454_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_2405_ _2408_/A _2405_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3842__B _3830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_221 VGND VPWR sky130_fd_sc_hd__fill_2
X_3385_ _2905_/A _2877_/X _3332_/C _2872_/B _3385_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2739__A _2727_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_574 VGND VPWR sky130_fd_sc_hd__fill_2
X_2336_ _2337_/A _2336_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4436__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_118 VGND VPWR sky130_fd_sc_hd__decap_4
X_2267_ _2253_/A _2272_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4376__D _3652_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_298 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_419 VGND VPWR sky130_fd_sc_hd__decap_6
X_4006_ _3993_/B _4005_/X _2602_/X _4552_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_65_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_611 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2474__A _2472_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_2198_ _2199_/A _2198_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2905__C _2900_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4586__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_357 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4413__RESET_B _2399_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3289__B _3275_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2984__B1 _3451_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_473 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_602 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2640__C _2639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_15 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2649__A _4522_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_585 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_478 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4286__D _2537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3190__D _3165_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_408 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_641 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_611 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2384__A _2388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_441 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_357 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_699 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3199__B _3144_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3927__B _2585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_501 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3646__C _3498_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4104__A _4105_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2727__B1 _3657_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3943__A _3943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_649 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4459__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3662__B _3430_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2559__A _4489_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3152__B1 _3095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_202 VGND VPWR sky130_fd_sc_hd__fill_2
X_3170_ _3219_/A _3122_/Y _3171_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_120_181 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_533 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2709__D _3816_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_268 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_611 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2294__A _2288_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2725__C _2527_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_493 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_176 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_305 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_647 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2966__B1 _2965_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3837__B _3830_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2954_ _2917_/B _2954_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2885_ _4376_/Q _2896_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2741__B _2741_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4204__A2_N _2741_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_4555_ _4555_/D _4555_/Q _2229_/X _4619_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4183__A2 _4180_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3506_ _3506_/A _3513_/B _3507_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3853__A _4535_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_627 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_115 VGND VPWR sky130_fd_sc_hd__decap_3
X_4486_ _4486_/D _4486_/Q _2312_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3930__A2 _3927_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3437_ _3503_/A _3437_/B _3437_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2469__A _2472_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_3368_ _2851_/X _3365_/X _3367_/X _3368_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__3143__B1 _3142_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_693 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3694__B2 _3693_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2319_ _2318_/A _2319_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_533 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_192 VGND VPWR sky130_fd_sc_hd__fill_2
X_3299_ _3280_/X _3297_/X _3298_/X _3297_/A _3277_/X _3300_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_57_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_205 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_132 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_688 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2932__A _3289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_636 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2957__B1 _2900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4601__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_432 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_498 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_487 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3482__B _3479_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_435 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2379__A _2379_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_360 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_181 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_235 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_202 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_555 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_536 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4335__RESET_B _2492_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_655 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3988__A2 _3979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_463 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3003__A _3003_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_603 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2842__A inport_data_i[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_636 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__B _2763_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_207 VGND VPWR sky130_fd_sc_hd__fill_2
X_2670_ _2666_/X _2670_/B _2670_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3673__A _3673_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3373__B1 _3372_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4569__SET_B _2213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_636 VGND VPWR sky130_fd_sc_hd__decap_4
X_4340_ _3313_/Y _2986_/A _2486_/X _4430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3392__B _3391_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_457 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2289__A _2288_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4271_ _4265_/A _4271_/B _4271_/C _4271_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_4_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_500 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3125__B1 _3095_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3222_ _3148_/A _3208_/A _3224_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_3153_ _3153_/A _3150_/X _3151_/Y _3153_/D _3153_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_94_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_566 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_257 VGND VPWR sky130_fd_sc_hd__fill_1
X_3084_ _3084_/A _3085_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2651__A2 _4526_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_422 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_124 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2752__A _4278_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3986_ _2701_/A _3986_/B _4554_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3567__B _3582_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2937_ _2936_/X _2979_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_179 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2902__D _2902_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2868_ _4378_/Q _2876_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4607_ _4255_/Y _4242_/A _2168_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3583__A _3554_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2799_ _2799_/A _2796_/X _2799_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4538_ _4538_/D _4538_/Q _2249_/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3903__A2 _3897_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_4469_ _3678_/X _4469_/Q _2332_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2199__A _2199_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_500 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_511 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2927__A _2926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_330 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_696 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2890__A2 _2887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_227 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_238 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4564__D _4564_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_400 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4092__A1 _3947_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_614 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3758__A _3759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_591 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_411 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_636 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2662__A _2657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_455 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_106 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3477__B _3475_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3493__A _3504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3355__B1 _3366_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_262 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4587__RESET_B _2191_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4516__RESET_B _2276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_680 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3658__A1 _3244_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_533 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_544 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_514 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2556__B _4488_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_577 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4474__D _4474_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2881__A2 _2880_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3668__A _3668_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_411 VGND VPWR sky130_fd_sc_hd__decap_12
X_3840_ _2657_/X _3827_/X _3839_/X _3840_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__2572__A _2571_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3771_ _3727_/X _3770_/B _3770_/X _3771_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_118_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_662 VGND VPWR sky130_fd_sc_hd__fill_1
X_2722_ _2721_/X _2722_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_538 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_695 VGND VPWR sky130_fd_sc_hd__fill_2
X_2653_ _2653_/A _2652_/X _2654_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3346__B1 _3347_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2584_ _3944_/B _2585_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_444 VGND VPWR sky130_fd_sc_hd__decap_4
X_4323_ _2845_/X _4323_/Q _2506_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_477 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_455 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_287 VGND VPWR sky130_fd_sc_hd__decap_6
X_4254_ _3388_/A _4264_/B _4254_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2747__A _4502_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4185_ _4185_/A _4185_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3205_ _3031_/X _3360_/A _3205_/C _3204_/X _3205_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_95_672 VGND VPWR sky130_fd_sc_hd__decap_4
X_3136_ _3041_/X _3068_/X _3066_/A _3045_/X _3136_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4384__D _3642_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3067_ _4356_/Q _3016_/Y _3071_/A _4355_/Q _3067_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_70_528 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4074__A1 _4570_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3578__A _3581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3821__A1 _2660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_422 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2482__A _2496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4082__A2_N _4081_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3297__B _3275_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_105 VGND VPWR sky130_fd_sc_hd__fill_2
X_3969_ _4568_/Q _3969_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_12_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3888__A1 _4541_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4202__A _4185_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_593 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_582 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4020__A2_N _4019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4559__D _4001_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_298 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3760__B _3760_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2657__A _4521_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4301__A2 _4299_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_171 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2807__D _2806_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_333 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_506 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_569 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3488__A _3488_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_399 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2392__A _2391_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2823__C _2822_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_263 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_477 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3935__B _2585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_694 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4469__D _3678_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_606 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3951__A _3950_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4350__RESET_B _2474_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_650 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2567__A _2604_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_536 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_366 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_528 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_26_0_clk_i_A clkbuf_4_13_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3398__A _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3823_ utmi_rxactive_i _3824_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_285 VGND VPWR sky130_fd_sc_hd__decap_3
X_3754_ _3745_/Y _3752_/X _3753_/Y _3754_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_118_346 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3845__B _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3685_ _4522_/Q _3685_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2705_ _2705_/A _2705_/B _2910_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_106_508 VGND VPWR sky130_fd_sc_hd__fill_2
X_2636_ _2636_/A _3707_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4438__RESET_B _2369_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4022__A _4564_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4379__D _4379_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_552 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3861__A _4538_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_19 VGND VPWR sky130_fd_sc_hd__fill_2
X_2567_ _2604_/A _2580_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2498_ _2497_/A _2498_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_436 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_414 VGND VPWR sky130_fd_sc_hd__fill_2
X_4306_ _2689_/B _3804_/B _2778_/X _4306_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3580__B _3583_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_257 VGND VPWR sky130_fd_sc_hd__decap_6
X_4237_ _4612_/Q _4237_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2477__A _2475_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_47 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_160 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2908__C _2908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4295__A1 _2524_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2845__A2 _2829_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4168_ _4168_/A _4188_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_28_558 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_355 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_344 VGND VPWR sky130_fd_sc_hd__fill_2
X_4099_ _4009_/X _4099_/B _4105_/A VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_15_208 VGND VPWR sky130_fd_sc_hd__decap_3
X_3119_ _3119_/A _3115_/X _3117_/X _3118_/X _3119_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4047__A1 _4565_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2924__B _2951_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_369 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_241 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3101__A _3221_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_285 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2940__A _3306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_469 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_99 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3474__C _3473_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4342__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_646 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_574 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_425 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3490__B _3488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2387__A _2388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4492__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_300 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3089__A2 _3088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_480 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2537__D _3820_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2834__B inport_accept_o VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3649__C _3648_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3797__B1 _2645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_591 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3011__A _4358_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2850__A _2905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3665__B _2826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4531__RESET_B _2258_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2772__B2 _2765_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3384__C _3384_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3470_ _3486_/B _3478_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_495 VGND VPWR sky130_fd_sc_hd__fill_2
X_2421_ _2419_/A _2421_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3316__A3 _3315_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_500 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3721__B1 _2673_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_2352_ _2352_/A _2352_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_3 VGND VPWR sky130_fd_sc_hd__decap_6
X_2283_ _2283_/A _2283_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2297__A _2301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_690 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_577 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_4022_ _4564_/Q _4022_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_439 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_620 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2827__A2 _2796_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_612 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_377 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3788__B1 _4488_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4017__A utmi_data_out_o[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3856__A _4536_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_611 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4365__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3806_ _3806_/A _3805_/X _3806_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4619__RESET_B _2155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2760__A _4497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3004__A2 _3003_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3136__A2_N _3068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_255 VGND VPWR sky130_fd_sc_hd__fill_2
X_3737_ _3724_/A _3737_/B _3736_/X _3737_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3575__B _3573_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_47 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_187 VGND VPWR sky130_fd_sc_hd__fill_2
X_3668_ _3668_/A _3668_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_109_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_29 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3591__A _3587_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3599_ _3585_/X _3597_/X _3598_/X _3599_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_2619_ _2618_/X _2796_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3712__B1 _3704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_555 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_266 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_22 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_333 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2935__A _2934_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2960__A2_N _3257_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2654__B _2654_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_472 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_686 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_174 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3779__B1 _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_122 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4572__D _4086_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3469__C _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_701 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3794__A3 _4490_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_76 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3188__D _3188_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_723 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3766__A _3762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2670__A _2666_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_255 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3485__B _3478_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_288 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_299 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_clk_i clkbuf_3_7_0_clk_i/A clkbuf_3_7_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__2754__A1 _2548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_509 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_454 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3703__B1 _3720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_406 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3006__A _3005_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2809__A2 _2784_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_322 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_50 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_333 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4482__D _3761_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_196 VGND VPWR sky130_fd_sc_hd__fill_2
X_2970_ _3491_/A _2969_/X _3491_/A _2969_/X _2970_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__4388__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_391 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_594 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3676__A _3669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2580__A _2580_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_597 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2730__D _2730_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4571_ _4571_/D _3931_/A _2211_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3522_ _3522_/A _3516_/B _3523_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3942__B1 _2552_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_658 VGND VPWR sky130_fd_sc_hd__decap_6
X_3453_ _3516_/A _3462_/B _3453_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2404_ _2408_/A _2404_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3384_ _3397_/A _3380_/X _3384_/C _4361_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_84_203 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_9_0_clk_i clkbuf_5_9_0_clk_i/A _4450_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_2335_ _2337_/A _2335_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_597 VGND VPWR sky130_fd_sc_hd__fill_1
X_2266_ _2261_/A _2266_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_428 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_247 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_642 VGND VPWR sky130_fd_sc_hd__decap_4
X_2197_ _2199_/A _2197_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4005_ _3994_/A _4552_/Q _4005_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_25_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_15 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4392__D _4392_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_431 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2681__B1 _2680_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2905__D _2904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3586__A _3498_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2984__B2 _3303_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4453__RESET_B _2351_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2490__A _2495_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_564 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_124 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_12 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4210__A _2706_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_553 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_435 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_446 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4567__D _4055_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_620 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2665__A _2671_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4110__B1 _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4530__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_306 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3496__A _3504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_513 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3646__D _3528_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2727__A1 outport_accept_i VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4104__B _4103_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3924__B1 _2610_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_317 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3662__C _3661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4120__A _2579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_691 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_680 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4477__D _3732_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2559__B _4488_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3152__A1 _3088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_545 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_193 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4101__B1 _3957_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2575__A _2575_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_461 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_601 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_196 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2725__D _2525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_144 VGND VPWR sky130_fd_sc_hd__decap_8
X_2953_ _2900_/D _3265_/B _2900_/D _3265_/B _2953_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_62_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_328 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2966__A1 _4331_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2884_ _2872_/B _2875_/X _2883_/X _2884_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__2741__C _2716_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_422 VGND VPWR sky130_fd_sc_hd__fill_2
X_4554_ _4554_/D _4554_/Q _2230_/X _4619_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3505_ _4411_/Q _3512_/B _3505_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4403__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3853__B _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_488 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_477 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_606 VGND VPWR sky130_fd_sc_hd__decap_6
X_4485_ _3779_/X _3674_/D _2313_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_89_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4030__A _4029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3930__A3 _3928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_127 VGND VPWR sky130_fd_sc_hd__fill_2
X_3436_ _3431_/X _3437_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3143__A1 _3029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_37 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4387__D _4387_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3367_ _3367_/A _3367_/B _3367_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_2318_ _2318_/A _2318_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4553__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3298_ _3253_/A _3298_/B _3298_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2485__A _2485_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2249_ _2248_/A _2249_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_420 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_250 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_12 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_114 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_199 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2957__B2 _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2932__B _2972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_372 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4205__A _2706_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_411 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_538 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_447 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_650 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_534 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2395__A _2391_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_431 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_623 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4375__RESET_B _2444_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3003__B _3248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_103 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_84 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2842__B _2846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_136 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__C _3656_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4426__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_387 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3373__A1 _2851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_560 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4576__CLK _4574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_447 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_4270_ _4270_/A _4264_/B _4271_/C VGND VPWR sky130_fd_sc_hd__nor2_4
X_3221_ _3221_/A _3112_/A _3218_/X _3220_/X _3221_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3125__A1 _3019_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_214 VGND VPWR sky130_fd_sc_hd__fill_2
X_3152_ _3088_/Y _3080_/Y _3095_/X _3153_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_67_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4086__C1 _4085_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3083_ _3082_/X _3084_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_82_559 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_637 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2752__B _2761_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3985_ _3984_/Y _3979_/X _3921_/Y _3981_/X _3986_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_2936_ _3297_/A _2935_/X _2936_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_50_478 VGND VPWR sky130_fd_sc_hd__fill_2
X_2867_ _2867_/A _4403_/Q _2862_/X _2866_/X _2867_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_109_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_208 VGND VPWR sky130_fd_sc_hd__fill_2
X_4606_ _4247_/X _4249_/A _2169_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3583__B _3583_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2798_ _2694_/A _2692_/Y _2633_/B _2799_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_7_90 VGND VPWR sky130_fd_sc_hd__decap_4
X_4537_ _4537_/D _4537_/Q _2250_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_296 VGND VPWR sky130_fd_sc_hd__fill_2
X_4468_ _2826_/X _4468_/Q _2333_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_89_169 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_147 VGND VPWR sky130_fd_sc_hd__fill_2
X_3419_ _3419_/A _3528_/B _3420_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_4399_ _4399_/D _2855_/A _2415_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_98_681 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_642 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_631 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2875__B1 _2874_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_567 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_526 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_6_0_clk_i clkbuf_4_7_0_clk_i/A clkbuf_4_6_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_589 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3104__A _3103_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_397 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_420 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4092__A2 _4056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3758__B _3770_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_261 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4575__SET_B _2205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_626 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_497 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2662__B _2658_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__CLK _4450_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4580__D _4147_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_158 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3477__C _3477_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_21 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4599__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__B _3491_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3355__A1 _3352_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_357 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_296 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_117 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3658__A2 _3657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_504 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2556__C _4486_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4556__RESET_B _2228_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3014__A _3013_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4068__C1 _4067_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2853__A _3634_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3949__A _4565_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_592 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3291__B1 _3289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_423 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4490__D _3794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_456 VGND VPWR sky130_fd_sc_hd__fill_2
X_3770_ _3727_/X _3770_/B _3770_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_630 VGND VPWR sky130_fd_sc_hd__fill_2
X_2721_ _2720_/X _2721_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_2652_ _2646_/Y _2647_/Y _2648_/X _2651_/X _2652_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_66_3 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3346__A1 _3347_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2583_ _2557_/X _3944_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_200 VGND VPWR sky130_fd_sc_hd__fill_1
X_4322_ _4322_/D _4322_/Q _2507_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4253_ _4253_/A _4264_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_489 VGND VPWR sky130_fd_sc_hd__decap_8
X_3204_ _3065_/X _3122_/Y _3204_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_95_640 VGND VPWR sky130_fd_sc_hd__decap_12
X_4184_ _4201_/A _4183_/X _4184_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_67_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_353 VGND VPWR sky130_fd_sc_hd__fill_2
X_3135_ _3055_/X _3098_/Y _3207_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_103_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_397 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_386 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2609__B1 _2608_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3066_ _3066_/A _3065_/X _3205_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3859__A _4537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2763__A _2763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4074__A2 _4056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_389 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3821__A2 _3804_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_283 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3578__B _3576_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_456 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3968_ _3967_/X utmi_data_out_o[6] VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_23_489 VGND VPWR sky130_fd_sc_hd__decap_6
X_2919_ _2918_/X _2920_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_3899_ _4546_/Q _3897_/X _3898_/X _3899_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3594__A _2857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_305 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4202__B _4194_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3888__A2 _3883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_629 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2938__A _3302_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_0_0_clk_i_A clkbuf_5_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3760__C _3759_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_331 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_320 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4575__D _4107_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_718 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_209 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2673__A _4520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_412 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3488__B _3478_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_445 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_622 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_143 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3009__A _4359_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_176 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_117 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2848__A inport_valid_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2839__B1 _2838_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4485__D _3779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4390__RESET_B _2427_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_301 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4614__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_60 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_526 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3679__A _3679_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_82 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_345 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_378 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2583__A _2557_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_721 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_272 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3398__B _3398_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_231 VGND VPWR sky130_fd_sc_hd__decap_6
X_3822_ _3822_/A _3822_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_60_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_415 VGND VPWR sky130_fd_sc_hd__fill_1
X_3753_ _3745_/Y _3752_/X _3720_/A _3753_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_9_460 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_3684_ _2660_/X _3669_/C _2660_/X _3669_/C _3684_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_493 VGND VPWR sky130_fd_sc_hd__fill_2
X_2704_ _2704_/A _2706_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2635_ _2635_/A _2636_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3861__B _3859_/B VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0_clk_i clkbuf_0_clk_i/X clkbuf_2_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4305_ _4467_/Q _2782_/X _4304_/X _4305_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_2566_ _2565_/X _2566_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2497_ _2497_/A _2497_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4407__RESET_B _2406_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_225 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_297 VGND VPWR sky130_fd_sc_hd__fill_2
X_4236_ _4236_/A _4236_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_59_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_26 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4395__D _3565_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2908__D _2907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4295__A2 _2725_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4167_ _4197_/A _4167_/B _4166_/Y _4585_/D VGND VPWR sky130_fd_sc_hd__and3_4
X_3118_ _3098_/Y _3094_/X _3219_/A _3118_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_83_676 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3589__A _3610_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_367 VGND VPWR sky130_fd_sc_hd__decap_4
X_4098_ _3955_/A _4039_/B _4033_/A _4097_/X _4098_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4047__A2 _4037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3255__B1 _2917_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2493__A _2495_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_581 VGND VPWR sky130_fd_sc_hd__fill_2
X_3049_ _3350_/C _3016_/Y _4354_/Q _3120_/B _3049_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_82_197 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_562 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3101__B _3171_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_448 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_45 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_303 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2940__B _2940_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_38 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4213__A _2711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_531 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4235__A1_N _4234_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2668__A _2667_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3490__C _3490_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_662 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_651 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_312 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_548 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3499__A _3498_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_clk_i clkbuf_3_3_0_clk_i/A clkbuf_4_7_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_74_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_345 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_315 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3797__B2 _3792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3797__A1 _2601_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_551 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_306 VGND VPWR sky130_fd_sc_hd__decap_6
X_2420_ _2419_/A _2420_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3962__A _4559_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3721__B2 _3674_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3721__A1 _2643_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_713 VGND VPWR sky130_fd_sc_hd__fill_2
X_2351_ _2352_/A _2351_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4081__A2_N _4566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2578__A _3925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_523 VGND VPWR sky130_fd_sc_hd__decap_12
X_2282_ _2283_/A _2282_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4500__RESET_B _2294_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_589 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_109 VGND VPWR sky130_fd_sc_hd__decap_12
X_4021_ _4015_/X _4020_/X _4015_/X _4020_/X _4099_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_315 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3788__B2 _3786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3788__A1 _2657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3202__A _3137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_370 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3856__B _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3805_ _3804_/Y _3805_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2760__B _2730_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_5_0_clk_i clkbuf_5_4_0_clk_i/A _4574_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_3736_ _3736_/A _3734_/X _3736_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3575__C _3574_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4033__A _4033_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_267 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3872__A _3824_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3667_ _3667_/A _3683_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4479__SET_B _2320_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3598_ outport_data_o[2] _3592_/B _3598_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2618_ _4514_/Q _2784_/A _2618_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3712__A1 _3708_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_512 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2488__A _2485_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2549_ _2519_/Y _2547_/X _4468_/Q _2548_/Y _2549_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_114_383 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_278 VGND VPWR sky130_fd_sc_hd__decap_12
X_4219_ _4219_/A _2548_/Y _4469_/Q _4219_/D _4219_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_28_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_67 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_78 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3779__A1 _3724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_11 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3112__A _3112_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3469__D _3528_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2951__A _2951_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_212 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3766__B _3764_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2670__B _2670_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3400__B1 _3412_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_216 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2754__A2 _4282_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_249 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_188 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3782__A _3785_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_400 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4329__RESET_B _2499_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3703__A1 _3702_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2398__A _2399_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_372 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_702 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_223 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_74 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_364 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_267 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_109 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3006__B _3216_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_632 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4118__A _4115_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3022__A _4355_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3957__A _4566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2861__A _2860_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_573 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_584 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3676__B _3672_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4570_ _4570_/D _4570_/Q _2212_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3521_ _2866_/A _3513_/B _3521_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3942__A1 _2578_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_615 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3942__B2 _3941_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3452_ outport_data_o[4] _3516_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2403_ _2396_/A _2408_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_201 VGND VPWR sky130_fd_sc_hd__decap_4
X_3383_ _3366_/A _3381_/X _3383_/C _3384_/C VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_111_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_212 VGND VPWR sky130_fd_sc_hd__fill_2
X_2334_ _2337_/A _2334_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_245 VGND VPWR sky130_fd_sc_hd__decap_6
X_2265_ _2261_/A _2265_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_2196_ _2199_/A _2196_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4004_ _2736_/X _4003_/X _4560_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_53_624 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4028__A _4562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_315 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4332__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2681__A1 _3780_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_635 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3867__A _4541_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_465 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_28_0_clk_i clkbuf_5_29_0_clk_i/A _4418_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_52_178 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_510 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4482__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3586__B _3528_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_486 VGND VPWR sky130_fd_sc_hd__fill_2
X_3719_ _3704_/A _3719_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4493__RESET_B _2304_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_7 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4422__RESET_B _2388_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4210__B _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3697__B1 _3684_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3107__A _3068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_458 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_237 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2665__B _2631_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4110__B2 _4562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_451 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_10 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4583__D _4583_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_646 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_476 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_679 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_498 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3496__B _3494_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_565 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2727__A2 _2725_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3924__A1 _2610_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3924__B2 _3923_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_263 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3688__B1 _2674_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2559__C _2522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4120__B _2572_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3152__A2 _3080_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3017__A _3015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_576 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_684 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_513 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2856__A _4397_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_72 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_61 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4355__CLK _4356_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_557 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4101__A1 _4566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4101__B2 _3966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2575__B _4437_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4493__D _3797_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_473 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_624 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3860__B1 _3859_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_410 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_635 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_clk_i clkbuf_2_1_0_clk_i/A clkbuf_2_0_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_50_605 VGND VPWR sky130_fd_sc_hd__decap_4
X_2952_ _4330_/Q _2922_/B _2951_/Y _3265_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3687__A _3687_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2591__A _2591_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_381 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2966__A2 _2951_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2883_ _2881_/Y _2882_/X _2883_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2741__D _2740_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_373 VGND VPWR sky130_fd_sc_hd__decap_8
X_4553_ _4553_/D _4553_/Q _2232_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3504_ _3504_/A _3504_/B _3504_/C _4410_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_116_445 VGND VPWR sky130_fd_sc_hd__fill_2
X_4484_ _3775_/X _3673_/A _2314_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_7_580 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_467 VGND VPWR sky130_fd_sc_hd__fill_2
X_3435_ outport_data_o[0] _3503_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_3366_ _3366_/A _3343_/Y _3367_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3143__A2 _3061_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2317_ _2324_/A _2318_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_384 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2974__A2_N _2973_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2766__A _4491_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3297_ _3297_/A _3275_/B _3297_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2248_ _2248_/A _2248_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_122_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_590 VGND VPWR sky130_fd_sc_hd__decap_3
X_2179_ _2177_/A _2179_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_25_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_668 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3597__A _2859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_498 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_24 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_295 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_690 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4205__B _2754_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4603__RESET_B _2172_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk_i clkbuf_4_3_0_clk_i/A clkbuf_5_4_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_119_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_456 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_467 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4578__D _4129_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4378__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_211 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2676__A _2675_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_505 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_97 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_495 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_81 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_498 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3300__A _3279_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__D _3657_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_195 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4344__RESET_B _2481_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3373__A2 _3370_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4131__A _2562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4488__D _3788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3970__A _4324_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_82 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3125__A2 _3026_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3220_ _3108_/X _3137_/A _3220_/C _3219_/X _3220_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_79_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_524 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2586__A _2560_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3074__A2_N _3070_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3151_ _3046_/X _3008_/X _3369_/A _3151_/D _3151_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_39_226 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_579 VGND VPWR sky130_fd_sc_hd__fill_2
X_3082_ _4358_/Q _4359_/Q _3007_/X _3008_/X _3082_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4086__B1 _4050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3833__B1 _3832_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_251 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4306__A _2689_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_402 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_446 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3210__A _4348_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_137 VGND VPWR sky130_fd_sc_hd__decap_12
X_3984_ _3984_/A _3984_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2935_ _2934_/X _2935_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2866_ _2866_/A _2863_/X _2864_/X _2865_/X _2866_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_4605_ _4605_/D _3413_/A _2170_/X _4619_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2797_ _2788_/A _2796_/X _4508_/Q _2797_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__4010__B1 _4008_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4041__A _4041_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4536_ _3876_/X _4536_/Q _2251_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4398__D _3575_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4520__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_48 VGND VPWR sky130_fd_sc_hd__fill_2
X_4467_ _4305_/X _4467_/Q _2334_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_104_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_4398_ _3575_/Y _2855_/B _2416_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3418_ _3427_/B _3528_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_77_19 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_0_0_clk_i_A clkbuf_4_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2496__A _2496_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3349_ _3397_/A _3345_/X _3349_/C _3349_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_112_492 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_343 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2875__A1 _2861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_605 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_273 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2662__C _2653_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_446 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4216__A _2750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3120__A _3071_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_660 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_693 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3493__C _3493_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3355__A2 _3354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_286 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3790__A _2669_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_418 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_693 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_365 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_354 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4068__B1 _4050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_324 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_549 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3815__B1 _3814_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2556__D _2523_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_432 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_571 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3291__B2 _3277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3291__A1 _3280_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2853__B _3643_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_476 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4596__RESET_B _2180_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_402 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4525__RESET_B _2265_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3030__A _3029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_435 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_619 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4543__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2720_ _2715_/X _4278_/D _2720_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_130 VGND VPWR sky130_fd_sc_hd__decap_3
X_2651_ _2649_/Y _4526_/Q _4522_/Q _2650_/Y _2651_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_8_185 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3346__A2 _3325_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2582_ _2581_/X _4552_/Q _2582_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_113_223 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3751__C1 _3750_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4321_ _2841_/X _4321_/Q _2508_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_608 VGND VPWR sky130_fd_sc_hd__fill_2
X_4252_ _4242_/Y _4263_/B _4252_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_86_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_3203_ _2996_/A _3195_/Y _3203_/C _3203_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_95_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_4183_ _4182_/Y _4180_/Y _4182_/A _4180_/A _4183_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3205__A _3031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_140 VGND VPWR sky130_fd_sc_hd__decap_12
X_3134_ _3176_/A _3088_/Y _3137_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_538 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2609__A1 _2605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_229 VGND VPWR sky130_fd_sc_hd__fill_2
X_3065_ _3039_/Y _3369_/A _3046_/X _3375_/A _3065_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__3859__B _3859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_357 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2944__A1_N _3455_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_571 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2763__B _2763_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3578__C _3578_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_593 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_232 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4036__A _4030_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_446 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_3967_ _2579_/X _3965_/X _2552_/X _3966_/Y _3967_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_23_479 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3875__A _4544_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2918_ _4328_/Q _2918_/B _2918_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_10_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_3898_ utmi_data_in_i[2] _3895_/B _3898_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2793__B1 _2791_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3594__B _3589_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2849_ _2849_/A _2905_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4202__C _4198_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4519_ _4519_/D _4519_/Q _2272_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_713 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2938__B _2979_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4298__B1 _4297_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4416__CLK _4410_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_685 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_376 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_484 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2954__A _2917_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_324 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_4_0_clk_i_A clkbuf_5_4_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_10 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_402 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4591__D _4197_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_593 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4566__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3785__A _3785_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_100 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_540 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_667 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_656 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4289__B1 _2533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2848__B _2829_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2839__A1 _4320_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3025__A _3016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2864__A _4410_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_72 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_530 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_593 VGND VPWR sky130_fd_sc_hd__fill_1
X_3821_ _2660_/X _3804_/B _3820_/X _3821_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_60_552 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_265 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3695__A _3695_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_315 VGND VPWR sky130_fd_sc_hd__decap_6
X_3752_ _3683_/Y _3690_/A _3683_/A _3690_/Y _3752_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2775__B1 _4266_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_3683_ _3683_/A _3683_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_472 VGND VPWR sky130_fd_sc_hd__decap_8
X_2703_ _2702_/X _2704_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_2634_ _4516_/Q _2635_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2565_ _4620_/D _3994_/A _2565_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_221 VGND VPWR sky130_fd_sc_hd__fill_2
X_4304_ _2639_/X _2800_/X _2815_/X _2824_/X _4304_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_99_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_2496_ _2496_/A _2497_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_59_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4439__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4235_ _4234_/Y _4368_/Q _4232_/Y _4257_/A _4235_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4166_ _4164_/Y _4163_/C _4166_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
Xclkbuf_5_1_0_clk_i clkbuf_5_1_0_clk_i/A _4596_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_95_493 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_685 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_173 VGND VPWR sky130_fd_sc_hd__decap_6
X_3117_ _3347_/A _3035_/X _3014_/Y _3117_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_28_527 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_195 VGND VPWR sky130_fd_sc_hd__fill_2
X_4097_ _4093_/X _4095_/X _4096_/Y _4097_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4589__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3255__A1 _3251_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3255__B2 _3248_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_571 VGND VPWR sky130_fd_sc_hd__decap_4
X_3048_ _3047_/X _3048_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_70_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4204__B1 _2718_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_326 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2518__B1 _2763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_554 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_543 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4586__D _4171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_140 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_633 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_173 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2684__A _2669_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3797__A2 _3785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_585 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3706__C1 _3705_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2859__A _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3721__A2 _3673_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2350_ _2352_/A _2350_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_535 VGND VPWR sky130_fd_sc_hd__decap_6
X_2281_ _2253_/A _2283_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4496__D _4496_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_408 VGND VPWR sky130_fd_sc_hd__fill_2
X_4020_ _4016_/Y _4019_/X _4016_/Y _4019_/X _4020_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_324 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4540__RESET_B _2247_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_644 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_143 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_132 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_335 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2594__A _4050_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3788__A2 _3782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3202__B _3202_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_574 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4314__A enable_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_602 VGND VPWR sky130_fd_sc_hd__fill_2
X_3804_ _2601_/A _3804_/B _3804_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_118_112 VGND VPWR sky130_fd_sc_hd__fill_1
X_3735_ _3736_/A _3734_/X _3737_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_118_145 VGND VPWR sky130_fd_sc_hd__decap_4
X_3666_ _2826_/X _3677_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_3597_ _2859_/B _3589_/X _3597_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2769__A _4240_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3173__B1 _3095_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2617_ _2595_/A _4033_/A _2516_/X _2616_/X _2617_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3712__A2 _4472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_2548_ _2548_/A _2548_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_114_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_535 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_24_0_clk_i clkbuf_5_25_0_clk_i/A _4534_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4218_ _4281_/A _2546_/B _2733_/A _4219_/D VGND VPWR sky130_fd_sc_hd__o21a_4
X_2479_ _2475_/X _2479_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_493 VGND VPWR sky130_fd_sc_hd__decap_4
X_4149_ _4153_/A _4147_/C _4151_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_346 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_677 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3779__A2 _3674_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_135 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3112__B _3112_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2987__B1 _2986_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_563 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_371 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_56 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4224__A _2753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_707 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_123 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3400__A1 _3399_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_11 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4604__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_228 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_44 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_12_0_clk_i_A clkbuf_4_6_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2679__A _2657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2775__A1_N _4236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_434 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3703__A2 _3701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_478 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4369__RESET_B _2451_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_257 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_493 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3303__A _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_614 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4118__B _4116_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4485__SET_B _2313_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3676__C _3676_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4134__A _2736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3520_ _3514_/A _3518_/Y _3520_/C _4415_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_115_104 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3942__A2 _3940_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_649 VGND VPWR sky130_fd_sc_hd__decap_3
X_3451_ _3451_/A _3434_/B _3451_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_6_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2589__A _2579_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2402_ _2399_/A _2402_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_41_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_3382_ _3382_/A _3376_/Y _3383_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3155__B1 _3088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_235 VGND VPWR sky130_fd_sc_hd__fill_2
X_2333_ _2337_/A _2333_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_332 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_2264_ _2261_/A _2264_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_611 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4309__A _2159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_2195_ _2166_/X _2199_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4003_ _4002_/Y _3994_/B _3972_/Y _3981_/X _4003_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_65_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_603 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_71 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2681__A2 _2629_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4028__B _4027_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_39 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2969__B1 _2968_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3867__B _3859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_382 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_522 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3586__C _3498_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_443 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3883__A _3883_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3718_ _3708_/X _3683_/A _3704_/X _3717_/X _3718_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__2499__A _2497_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3649_ _3581_/A _3649_/B _3648_/X _3649_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_0_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3697__B2 _3696_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_170 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3107__B _3151_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_566 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4462__RESET_B _2341_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_365 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_600 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4219__A _4219_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_644 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2665__C _2664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_455 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_135 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_319 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3496__C _3495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_599 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3924__A2 _3922_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_500 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2202__A _2166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_253 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3688__A1 _4524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3688__B2 _2658_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2559__D _2525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_286 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4120__C _2575_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3017__B _3016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_544 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2856__B _3566_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_588 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_238 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_290 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4101__A2 _4007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4129__A _2736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2575__C _2575_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3033__A _4357_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3860__A1 _4529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_485 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3968__A _3967_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2872__A _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_2951_ _2951_/A _2951_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2591__B _2577_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_308 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_2882_ _2878_/Y _2861_/X _2880_/A _2879_/X _2882_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_4552_ _4552_/D _4552_/Q _2233_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3503_ _3503_/A _3513_/B _3504_/C VGND VPWR sky130_fd_sc_hd__and2_4
X_4483_ _3768_/X _3674_/B _2315_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_116_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_319 VGND VPWR sky130_fd_sc_hd__decap_12
X_3434_ _2902_/D _3434_/B _3434_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3208__A _3208_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_i_A clkbuf_2_0_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_17 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_352 VGND VPWR sky130_fd_sc_hd__decap_8
X_3365_ _3039_/Y _3364_/B _3369_/B _3365_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_111_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_2316_ _2314_/A _2316_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_514 VGND VPWR sky130_fd_sc_hd__fill_2
X_3296_ _3279_/A _3295_/Y _3296_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_2247_ _2248_/A _2247_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_396 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_558 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_709 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4039__A _3923_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_441 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_260 VGND VPWR sky130_fd_sc_hd__decap_12
X_2178_ _2177_/A _2178_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2782__A _2781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_466 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3597__B _3589_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_477 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_680 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_262 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4111__A1_N _4026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_416 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4594__D _4204_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_43 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4095__A1 _3966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_591 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_647 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2692__A _2620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_628 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_152 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3300__B _3300_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_185 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_341 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3358__B1 _2907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_378 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_8 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4131__B _4130_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4384__RESET_B _2434_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4322__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3028__A _3015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_416 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3970__B _3960_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2867__A _2867_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_385 VGND VPWR sky130_fd_sc_hd__fill_2
X_3150_ _3021_/X _3105_/D _3350_/C _3150_/D _3150_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_121_493 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4472__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3081_ _3055_/X _3080_/Y _3148_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4086__A1 _3939_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3698__A _3698_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3833__A1 _4517_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_466 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_433 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_414 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4306__B _3804_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3983_ _2701_/A _3983_/B _4553_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_16_691 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_149 VGND VPWR sky130_fd_sc_hd__decap_4
X_2934_ _3293_/A _2933_/X _2934_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_672 VGND VPWR sky130_fd_sc_hd__fill_2
X_2865_ _3543_/A _2865_/B _2865_/C _4411_/Q _2865_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_31_683 VGND VPWR sky130_fd_sc_hd__fill_2
X_4604_ _4604_/D _2763_/B _2171_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4535_ _3874_/X _4535_/Q _2254_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2796_ _2796_/A _2796_/B _2793_/Y _2795_/Y _2796_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4010__B2 _4009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_243 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4041__B _4039_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_265 VGND VPWR sky130_fd_sc_hd__decap_8
X_4466_ _2783_/Y _2763_/C _2335_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4397_ _3571_/Y _4397_/Q _2418_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_89_138 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2777__A _2764_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3417_ _2763_/A _2763_/B _2763_/C _3417_/D _3427_/B VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_98_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_503 VGND VPWR sky130_fd_sc_hd__fill_2
X_3348_ _3346_/X _3347_/Y _3366_/A _3349_/C VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_85_311 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2875__A2 _2867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_clk_i_A clkbuf_4_5_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3279_ _3279_/A _3278_/Y _4332_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_85_388 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_591 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3401__A _3398_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2662__D _2661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_285 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4216__B _4216_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3120__B _3120_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4232__A _4608_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4345__CLK _4325_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4589__D _4184_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3764__A2_N _3763_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2687__A _3704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4495__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3790__B _3790_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_521 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_514 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_536 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_86 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_569 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4068__A1 _4569_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_314 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_528 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3815__A1 _2674_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_591 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_444 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2853__C _4384_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3291__A2 _3289_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3311__A _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_285 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_447 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_672 VGND VPWR sky130_fd_sc_hd__fill_2
X_2650_ _4526_/Q _2650_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_665 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4142__A _4135_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4499__D _3809_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_403 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3200__C1 _3199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3981__A _3980_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2581_ _2581_/A _2581_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3751__B1 _3719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2988__A2_N _2987_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4320_ _4320_/D _4320_/Q _2509_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_4_370 VGND VPWR sky130_fd_sc_hd__fill_2
X_4251_ _4253_/A _4263_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2597__A _3994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_279 VGND VPWR sky130_fd_sc_hd__fill_2
X_3202_ _3137_/X _3202_/B _3202_/C _3203_/C VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_79_193 VGND VPWR sky130_fd_sc_hd__fill_2
X_4182_ _4182_/A _4182_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3205__B _3360_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_664 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_344 VGND VPWR sky130_fd_sc_hd__fill_2
X_3133_ _2996_/A _3133_/B _3133_/C _3133_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_103_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_163 VGND VPWR sky130_fd_sc_hd__fill_1
X_3064_ _3038_/Y _3375_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2609__A2 _2577_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_369 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_583 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2763__C _2763_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_252 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3221__A _3221_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_425 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4368__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_266 VGND VPWR sky130_fd_sc_hd__fill_1
X_3966_ _4007_/A _3966_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_11_609 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3875__B _3877_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2917_ _2917_/A _2917_/B _2918_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_10_119 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_480 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_508 VGND VPWR sky130_fd_sc_hd__decap_12
X_3897_ _3883_/A _3897_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2793__B2 _2792_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2793__A1 _2636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4052__A utmi_data_out_o[0] VGND VPWR sky130_fd_sc_hd__diode_2
X_2848_ inport_valid_i _2829_/A _2848_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_541 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3891__A _3891_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_19 VGND VPWR sky130_fd_sc_hd__decap_12
X_2779_ _2778_/X _2779_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4202__D _4202_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_574 VGND VPWR sky130_fd_sc_hd__fill_2
X_4518_ _4518_/D _4518_/Q _2273_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3742__B1 _3741_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4449_ _2664_/X _4449_/Q _2356_/X _4450_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2300__A _2301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4298__A1 _3960_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_506 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_474 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_34 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_219 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_358 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4227__A _2601_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_230 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_5_8_0_clk_i_A clkbuf_5_9_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_561 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_241 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_255 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_19_0_clk_i clkbuf_4_9_0_clk_i/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_41_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_613 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_686 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_530 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_123 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3733__B1 _2641_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_74 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3306__A _3306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4289__A1 _4497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_362 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2210__A _2238_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_227 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2839__A2 _2831_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2864__B _4413_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_656 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_358 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4510__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_369 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_550 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4137__A _2628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3041__A _3040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_199 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_520 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2880__A _2880_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3820_ _3820_/A _3804_/Y _3820_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_60_542 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3976__A _2579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3695__B _3695_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3751_ _3726_/X _3711_/B _3719_/X _3750_/Y _3751_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__2775__B2 _4494_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_480 VGND VPWR sky130_fd_sc_hd__fill_2
X_2702_ _2595_/A _4050_/A _2702_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3682_ _3668_/X _3675_/B _3668_/X _3675_/B _3682_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_3 VGND VPWR sky130_fd_sc_hd__decap_6
X_2633_ _4514_/Q _2633_/B _2633_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_200 VGND VPWR sky130_fd_sc_hd__decap_6
X_2564_ _2705_/A _3994_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4303_ _4372_/Q _3420_/X _3660_/A _4303_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_87_428 VGND VPWR sky130_fd_sc_hd__decap_8
X_2495_ _2495_/A _2495_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3216__A _3216_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_288 VGND VPWR sky130_fd_sc_hd__fill_2
X_4234_ _4234_/A _4234_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_4_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_39 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_141 VGND VPWR sky130_fd_sc_hd__fill_2
X_4165_ _4164_/Y _4163_/C _4167_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_3116_ _3021_/X _3347_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4096_ _4093_/X _4095_/X _4030_/X _4096_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__3255__A2 _3253_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_701 VGND VPWR sky130_fd_sc_hd__fill_1
X_3047_ _3046_/X _3008_/X _3039_/Y _3010_/X _3047_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4487__RESET_B _2311_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_380 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_531 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_723 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3886__A _3824_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4416__RESET_B _2395_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2790__A _2694_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_233 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_586 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4204__B2 _4281_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_20_0_clk_i clkbuf_5_21_0_clk_i/A _4325_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3949_ _4565_/Q _3949_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_109_338 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3963__B1 _2581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_500 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2518__A1 _3416_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_393 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_115 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_566 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3126__A _3048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_11 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2965__A _2965_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4533__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_196 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2693__B1_N _2692_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3797__A3 _4493_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_520 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2205__A _2206_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3954__B1 _2604_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_432 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3706__B1 _3704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2859__B _2859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3036__A _3031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_547 VGND VPWR sky130_fd_sc_hd__fill_2
X_2280_ _2277_/A _2280_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_569 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_258 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_472 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_314 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_656 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_358 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_509 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_648 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3788__A3 _3790_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_328 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4580__RESET_B _2199_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3202__C _3202_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_572 VGND VPWR sky130_fd_sc_hd__decap_4
X_3803_ _3804_/B _3803_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_597 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_586 VGND VPWR sky130_fd_sc_hd__fill_2
X_3734_ _3679_/A _4472_/Q _3702_/A _3680_/Y _3734_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4406__CLK _4410_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3665_ _4469_/Q _2826_/X _3678_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_319 VGND VPWR sky130_fd_sc_hd__fill_2
X_2616_ utmi_txready_i _4029_/C _2591_/A _2616_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_114_330 VGND VPWR sky130_fd_sc_hd__decap_6
X_3596_ _3585_/X _3596_/B _3595_/X _4387_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_102_503 VGND VPWR sky130_fd_sc_hd__decap_6
X_2547_ _2520_/Y _2546_/X _2547_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3173__B2 _3122_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4556__CLK _4619_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2478_ _2475_/X _2478_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_547 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2785__A _2804_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4217_ _4214_/Y _4216_/X _4278_/D _4217_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_68_472 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_623 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_291 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_111 VGND VPWR sky130_fd_sc_hd__fill_2
X_4148_ _4581_/Q _4153_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_28_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_475 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_4079_ _4079_/A _4079_/B _4079_/C _4079_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_70_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_188 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3112__C _3190_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_158 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2987__A1 _2986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_383 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_715 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_575 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_719 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_102 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3400__A2 _3398_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_269 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_157 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4240__A _4240_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_691 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2679__B _2658_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4597__D _4209_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_311 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_396 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_16_0_clk_i_A clkbuf_4_8_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4113__B1 _4112_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_464 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3303__B _3303_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4338__RESET_B _2488_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_103 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4118__C _4117_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_74 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_512 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3676__D _3675_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4429__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4134__B _4132_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_589 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4579__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_138 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_116 VGND VPWR sky130_fd_sc_hd__fill_2
X_3450_ _3424_/X _3450_/B _3449_/X _3450_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA_clkbuf_2_0_0_clk_i_A clkbuf_2_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4150__A _4153_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3155__A1 _3219_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2589__B _2572_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2401_ _2399_/A _2401_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3381_ _3381_/A _3376_/A _3381_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_523 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_225 VGND VPWR sky130_fd_sc_hd__decap_3
X_2332_ _2337_/A _2332_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_3 VGND VPWR sky130_fd_sc_hd__decap_8
X_2263_ _2261_/A _2263_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_4002_ _4603_/Q _4002_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_84_239 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_133 VGND VPWR sky130_fd_sc_hd__decap_3
X_2194_ _2188_/X _2194_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_92_261 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_250 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_475 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_283 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_423 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2969__A1 _2926_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_681 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3586__D _3528_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_394 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_534 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_578 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_589 VGND VPWR sky130_fd_sc_hd__fill_2
X_3717_ _3717_/A _3674_/B _3717_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4040__C1 _4039_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_477 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_127 VGND VPWR sky130_fd_sc_hd__fill_2
X_3648_ _3547_/A _3646_/Y _3648_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4060__A _4061_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3579_ _4400_/Q _3582_/B _3579_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_416 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4219__B _2548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_79 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2665__D _2671_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_166 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4431__RESET_B _2377_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_34 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_199 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_78 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_670 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_361 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3909__B1 _3908_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_505 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_556 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_538 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_171 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3688__A2 _4525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_512 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_70 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_81 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3017__C _4354_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4519__RESET_B _2272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3314__A _3314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4098__C1 _4097_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4129__B _4119_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_604 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3860__A2 _3855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_648 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_199 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2872__B _2872_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_136 VGND VPWR sky130_fd_sc_hd__fill_2
X_2950_ _3494_/A _2949_/X _3494_/A _2949_/X _2950_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__2591__C utmi_txvalid_o VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4145__A _4146_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_361 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2820__B1 _2785_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2881_ _2878_/Y _2880_/X _2871_/B _2881_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4620_/D _3392_/A _4309_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3984__A _3984_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4551_ _3909_/X _3891_/A _2234_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_560 VGND VPWR sky130_fd_sc_hd__fill_2
X_3502_ _3516_/B _3513_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_4482_ _3761_/X _3715_/B _2316_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3433_ _3462_/B _3434_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3208__B _3176_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_331 VGND VPWR sky130_fd_sc_hd__fill_2
X_3364_ _3039_/Y _3364_/B _3369_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_686 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_2315_ _2314_/A _2315_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3295_ _3280_/X _3293_/X _3294_/X _3293_/A _3277_/X _3295_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_57_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4_0_clk_i_A clkbuf_2_2_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3224__A _3224_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2246_ _2248_/A _2246_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_537 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4564__SET_B _2219_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4039__B _4039_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_209 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_272 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_475 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_2177_ _2177_/A _2177_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2774__A1_N _4608_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2811__B1 _3704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_342 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_519 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2303__A _2324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_526 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4612__RESET_B _2161_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_11 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3134__A _3176_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4095__A2 utmi_data_out_o[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_423 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_61 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2692__B _2810_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_297 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_117 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_175 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_662 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_191 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3358__A1 _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_673 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_386 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3309__A _3317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2213__A _2210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4131__C _2587_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3028__B _3016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_406 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_106 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_40 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_574 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2867__B _4403_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4233__A1_N _4232_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_461 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4617__CLK _4619_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4353__RESET_B _2471_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3080_ _3079_/X _3080_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3044__A _3359_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4086__A2 _4056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3979__A _3994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3833__A2 _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_389 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2883__A _2881_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_670 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_618 VGND VPWR sky130_fd_sc_hd__fill_2
X_3982_ _4116_/A _3979_/X _3912_/Y _3981_/X _3983_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_90_595 VGND VPWR sky130_fd_sc_hd__decap_12
X_2933_ _2932_/X _2933_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4306__C _2778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11_0_clk_i_A clkbuf_3_5_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_2864_ _4410_/Q _4413_/Q _4412_/Q _2864_/D _2864_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_117_712 VGND VPWR sky130_fd_sc_hd__fill_2
X_2795_ _2624_/A _2654_/X _2794_/X _2795_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_4603_ _4603_/D _4603_/Q _2172_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4534_ _3871_/X _4534_/Q _2255_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3219__A _3219_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_255 VGND VPWR sky130_fd_sc_hd__decap_8
X_4465_ _4527_/Q outport_data_o[7] _2336_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4396_ _3568_/Y _3566_/A _2419_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2777__B _2767_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3416_ _3416_/A _4514_/Q _3419_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_85_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_515 VGND VPWR sky130_fd_sc_hd__decap_4
X_3347_ _3347_/A _3347_/B _3325_/X _3347_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3889__A _3889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_667 VGND VPWR sky130_fd_sc_hd__decap_12
X_3278_ _3251_/X _3275_/X _3276_/X _2926_/A _3277_/X _3278_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_85_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_581 VGND VPWR sky130_fd_sc_hd__decap_4
X_2229_ _2228_/A _2229_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_445 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_8_0_clk_i_A clkbuf_4_9_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3401__B _3400_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_618 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_595 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_297 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3120__C _3023_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_684 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_327 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3129__A _3129_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_222 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2968__A _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_29 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_15_0_clk_i clkbuf_4_7_0_clk_i/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_103_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_651 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_10 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_98 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4068__A2 _4056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3815__A2 _3803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_31 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3291__A3 _3290_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2853__D _2853_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3311__B _2987_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2208__A _2206_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_297 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_684 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4142__B _4137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3039__A _4358_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3200__B1 _3171_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2580_ _2580_/A _2581_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3751__A1 _3726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_415 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4534__RESET_B _2255_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2878__A _2877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_448 VGND VPWR sky130_fd_sc_hd__fill_1
X_4250_ _4249_/Y _4250_/B _4253_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_4181_ _4201_/A _4181_/B _4180_/Y _4181_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_3201_ _3209_/A _3198_/X _3200_/X _3202_/B VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_121_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_323 VGND VPWR sky130_fd_sc_hd__fill_2
X_3132_ _3132_/A _3129_/X _3202_/C _3133_/C VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_95_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3205__C _3205_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3267__B1 _4330_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_581 VGND VPWR sky130_fd_sc_hd__decap_3
X_3063_ _3010_/X _3369_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3502__A _3516_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_562 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2763__D _2725_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3221__B _3112_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4110__A1_N _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_392 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_275 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_256 VGND VPWR sky130_fd_sc_hd__fill_2
X_3965_ _2572_/X _3963_/Y _2611_/X _3964_/Y _3965_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3896_ _4545_/Q _3883_/X _3895_/X _3896_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_2916_ _2915_/X _2916_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_10_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2793__A2 _2790_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2847_ _4324_/Q _2829_/A _2846_/X _4324_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4052__B _4053_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3891__B _3895_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2778_ _2777_/X _2778_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_597 VGND VPWR sky130_fd_sc_hd__fill_1
X_4517_ _3833_/X _4517_/Q _2275_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3742__A1 _3680_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2788__A _2788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_225 VGND VPWR sky130_fd_sc_hd__fill_2
X_4448_ _4448_/D _2810_/B _2357_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4298__A2 _4292_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_632 VGND VPWR sky130_fd_sc_hd__decap_8
X_4379_ _4379_/D _4379_/Q _2440_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_665 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_710 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_721 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3412__A _3412_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_212 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_610 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4462__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_632 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_113 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3733__B2 _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2698__A _2654_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_718 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_707 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3306__B _3246_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4289__A2 _4286_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_654 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_643 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_30 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3249__B1 _2917_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_518 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2864__C _4412_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_646 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_713 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4137__B _4137_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2880__B _2879_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3976__B _3976_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3750_ _3708_/A _3748_/X _3749_/Y _3750_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4153__A _4153_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_429 VGND VPWR sky130_fd_sc_hd__fill_2
X_2701_ _2701_/A _2700_/Y _4448_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_118_328 VGND VPWR sky130_fd_sc_hd__fill_2
X_3681_ _3680_/Y _4474_/Q _3680_/Y _4474_/Q _3681_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3992__A _2701_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2632_ _2784_/A _2633_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_64_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_2563_ utmi_txready_i _2705_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2401__A _2399_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4302_ enable_i utmi_op_mode_o[0] VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_556 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_418 VGND VPWR sky130_fd_sc_hd__decap_8
X_2494_ _2495_/A _2494_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4233_ _4232_/Y _4257_/A _4612_/Q _3407_/Y _4233_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3216__B _3216_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_654 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_131 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_4164_ _4585_/Q _4164_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_315 VGND VPWR sky130_fd_sc_hd__decap_3
X_4095_ _3966_/Y utmi_data_out_o[7] _4094_/X _4095_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_3115_ _3061_/X _3018_/X _3094_/X _3114_/X _3115_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_82_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4335__CLK _4334_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3046_ _3007_/X _3046_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3763__A2_N _2660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3255__A3 _3254_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_178 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_551 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_189 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_201 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4485__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2790__B _2790_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3948_ _2571_/X _3946_/X _2611_/X _4046_/A _3948_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3963__A1 _2605_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3879_ _4546_/Q _3877_/B _3879_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_109_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4456__RESET_B _2348_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3963__B2 _3962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3701__A2_N _3700_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2518__A2 _4514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_628 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2311__A _2314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3407__A _4270_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_578 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_407 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3126__B _3150_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_526 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_304 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_186 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_337 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3142__A _3082_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_73 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_66 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_267 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3954__A1 _2581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3954__B2 _4558_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3706__A1 _3705_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_350 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_0_0_clk_i_A clkbuf_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_477 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2859__C _2859_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3317__A _3317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2221__A _2217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_418 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3036__B _3035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_515 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_215 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4358__CLK _4334_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_624 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4148__A _4581_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3890__B1 _3889_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2693__A1 _3720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3052__A _3048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_616 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_668 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3987__A _3987_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2891__A _2861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_595 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_543 VGND VPWR sky130_fd_sc_hd__decap_6
X_3802_ _3802_/A _3804_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_615 VGND VPWR sky130_fd_sc_hd__fill_1
X_3733_ _2641_/Y _3685_/X _2641_/Y _3685_/X _3736_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_259 VGND VPWR sky130_fd_sc_hd__decap_4
X_3664_ _3528_/A _3430_/A _3663_/X _3664_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_118_158 VGND VPWR sky130_fd_sc_hd__fill_2
X_2615_ utmi_txvalid_o _4029_/C VGND VPWR sky130_fd_sc_hd__inv_8
X_3595_ outport_data_o[1] _3592_/B _3595_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3227__A _3381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_2546_ _2724_/A _2546_/B _2546_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_2477_ _2475_/X _2477_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_237 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2785__B _4447_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4216_ _2750_/X _4216_/B _4216_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4147_ _4143_/X _4147_/B _4147_/C _4147_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_110_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_432 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_646 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_337 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3897__A _3883_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4078_ utmi_data_out_o[4] _4076_/X _4079_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_83_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3112__D _3111_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3029_ _3028_/X _3029_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2987__A2 _2986_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_340 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_587 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2306__A _2306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_114 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_670 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2679__C _2678_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4240__B _4240_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3137__A _3137_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_342 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_705 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4500__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_66 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_440 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4113__A1 _4109_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_218 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3321__C1 _3244_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_679 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_638 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3600__A _2859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_53 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4378__RESET_B _2441_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_351 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4134__C _4134_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_598 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2216__A _2210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_524 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2400_ _2399_/A _2400_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_109_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4150__B _4147_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2589__C _2582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3047__A _3046_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3380_ _3334_/X _3374_/X _3337_/Y _3380_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3155__A2 _3014_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_513 VGND VPWR sky130_fd_sc_hd__decap_4
X_2331_ _2324_/A _2337_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_2262_ _2261_/A _2262_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_4001_ _2736_/X _4000_/X _4001_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_77_292 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_646 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_123 VGND VPWR sky130_fd_sc_hd__decap_4
X_2193_ _2188_/X _2193_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_1_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_19 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_95 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3510__A _3510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2969__A2 _2965_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3733__A1_N _2641_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_170 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_546 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4040__B1 _4033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_423 VGND VPWR sky130_fd_sc_hd__decap_4
X_3716_ _3708_/X _4474_/Q _3704_/X _3715_/X _4474_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4523__CLK _4539_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_489 VGND VPWR sky130_fd_sc_hd__fill_2
X_3647_ _4375_/Q _3646_/Y _3649_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4060__B _4059_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3578_ _3581_/A _3576_/Y _3578_/C _4399_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_121_109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_513 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2796__A _2796_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2529_ _4615_/Q _4614_/Q _4616_/Q _2530_/C VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_0_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_389 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3854__B1 _3853_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_410 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4219__C _4469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_443 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_262 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_627 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3420__A _3420_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_446 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_52 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4400__RESET_B _2414_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3909__A1 _3891_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_56 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_517 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2957__A1_N _2900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4251__A _4253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_200 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4401__D _4401_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_524 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_31_0_clk_i_A clkbuf_5_30_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_20 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3017__D _4355_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_505 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4098__B1 _4033_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3314__B _3246_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_443 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4129__C _4128_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_91 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_413 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4559__RESET_B _2225_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3330__A _3327_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2872__C _2869_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4145__B _4137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4546__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2820__A1 _2636_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2880_ _2880_/A _2879_/X _2880_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_70_490 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_90 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_373 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4161__A _4187_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_398 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550_ _3907_/X _3889_/A _2235_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_550 VGND VPWR sky130_fd_sc_hd__decap_8
X_3501_ _4410_/Q _3512_/B _3504_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_116_426 VGND VPWR sky130_fd_sc_hd__fill_2
X_4481_ _4481_/D _3713_/B _2318_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_116_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_3432_ _3431_/X _3462_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3208__C _3206_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3363_ _3363_/A _3325_/X _3364_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3505__A _4411_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_665 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_376 VGND VPWR sky130_fd_sc_hd__fill_2
X_2314_ _2314_/A _2314_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3294_ _3243_/B _2946_/X _3294_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_207 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3836__B1 utmi_rxactive_i VGND VPWR sky130_fd_sc_hd__diode_2
X_2245_ _2238_/A _2248_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3224__B _3156_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2176_ _2177_/A _2176_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_605 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_104 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_616 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3240__A _3240_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_690 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_38 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2811__A1 _2699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_376 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4013__B1 utmi_data_out_o[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4071__A utmi_data_out_o[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_643 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3415__A _3508_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_654 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4419__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3134__B _3088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_508 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_432 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_627 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_476 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_498 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4246__A _4233_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_446 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4569__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3150__A _3021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_107 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_11_0_clk_i clkbuf_4_5_0_clk_i/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_685 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3358__A2 _3354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3309__B _3308_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4570__SET_B _2212_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_81 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4131__D _4118_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3028__C _3071_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2867__C _2862_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_52 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_343 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3325__A _3324_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_218 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3044__B _3043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4393__RESET_B _2422_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_560 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2883__B _2882_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_541 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4322__RESET_B _2507_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3060__A _3007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4156__A _4156_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4243__B1 _4236_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VPWR sky130_fd_sc_hd__decap_3
X_3981_ _3980_/X _3981_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2932_ _3289_/A _2972_/A _2932_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_62_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_2863_ _4414_/Q _2863_/B _2863_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2404__A _2408_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2794_ _2635_/A _2790_/B _2639_/X _2794_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4602_ _4602_/D _4602_/Q _2173_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_30_195 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_clk_i_A clkbuf_3_7_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4533_ _3868_/X _4533_/Q _2256_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3219__B _3026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_391 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_29 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_429 VGND VPWR sky130_fd_sc_hd__fill_2
X_4464_ _4526_/Q outport_data_o[6] _2337_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4395_ _3565_/Y _3563_/A _2420_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3415_ _3508_/A _3415_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2777__C _2768_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3346_ _3347_/A _3325_/X _3347_/B _3346_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_112_484 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3889__B _3895_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3277_ _3277_/A _3277_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3809__B1 _3808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_679 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_560 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_2228_ _2228_/A _2228_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_53_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_210 VGND VPWR sky130_fd_sc_hd__decap_12
X_2159_ _2159_/A _2163_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_284 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4066__A _4066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_424 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_449 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_438 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3120__D _3016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2314__A _2314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3129__B _3112_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3145__A _3079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_685 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4391__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_508 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_700 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_435 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_552 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4225__B1 _2745_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_601 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_634 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_482 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2224__A _2238_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3200__A1 _3045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4142__C _4197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3751__A2 _3711_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_394 VGND VPWR sky130_fd_sc_hd__decap_3
X_4180_ _4180_/A _4180_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3200_ _3045_/X _3014_/Y _3171_/B _3199_/Y _3200_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3055__A _3054_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_173 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2894__A _2893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3131_ _3085_/A _3066_/A _3130_/X _2997_/X _3202_/C VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_67_357 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4503__RESET_B _2291_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3205__D _3204_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3267__B2 _3248_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3267__A1 _3251_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_519 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_3062_ _3061_/X _3066_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_94_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_349 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_722 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3221__C _3218_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_224 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_298 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_287 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_246 VGND VPWR sky130_fd_sc_hd__decap_4
X_3964_ _3964_/A _3964_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3895_ utmi_data_in_i[1] _3895_/B _3895_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2915_ _3244_/B _3241_/A _2915_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2846_ inport_data_i[7] _2846_/B _2846_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2777_ _2764_/Y _2767_/X _2768_/Y _2776_/X _2777_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_117_565 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3742__A2 _3740_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4516_ _3831_/X _4516_/Q _2276_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_104_237 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_4447_ _4447_/D _4447_/Q _2358_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__2950__B1 _3494_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_611 VGND VPWR sky130_fd_sc_hd__fill_2
X_4378_ _3623_/X _4378_/Q _2441_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3329_ _4397_/Q _3566_/A _3329_/C _2855_/X _3329_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_58_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_390 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2309__A _2306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3412__B _3412_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_276 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_449 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4607__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3718__C1 _3717_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2979__A _2979_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_648 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_699 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2698__B _2662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_331 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_460 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_386 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_143 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3603__A _2858_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3249__B2 _3248_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3249__A1 _3243_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_700 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2864__D _2864_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_390 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_530 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_722 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2219__A _2217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_232 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_371 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_585 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_246 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4153__B _4153_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2700_ _4510_/Q _2810_/B _2687_/X _2699_/X _2700_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XFILLER_13_493 VGND VPWR sky130_fd_sc_hd__fill_2
X_3680_ _4472_/Q _3680_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3992__B _3991_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_486 VGND VPWR sky130_fd_sc_hd__fill_2
X_2631_ _2601_/A _3717_/A _2691_/A _2804_/A _2670_/B _2631_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__2889__A _3367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2562_ inport_valid_i _2557_/X _2908_/C _4278_/C _2562_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_114_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_213 VGND VPWR sky130_fd_sc_hd__fill_2
X_4301_ _4292_/Y _4299_/Y _4300_/Y _4619_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_114_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_2493_ _2495_/A _2493_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4232_ _4608_/Q _4232_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_4_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_590 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3513__A _3513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_19 VGND VPWR sky130_fd_sc_hd__fill_1
X_4163_ _4143_/X _4161_/Y _4163_/C _4163_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_82_102 VGND VPWR sky130_fd_sc_hd__fill_2
X_4094_ _3966_/Y utmi_data_out_o[7] _4094_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3114_ _3011_/X _3369_/A _3046_/X _3375_/A _3114_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_83_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_338 VGND VPWR sky130_fd_sc_hd__decap_4
X_3045_ _3044_/X _3045_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_82_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_596 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_408 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_419 VGND VPWR sky130_fd_sc_hd__fill_2
X_3947_ _3947_/A _4046_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_23_16 VGND VPWR sky130_fd_sc_hd__fill_2
X_3878_ _4537_/Q _3869_/X _3877_/X _4537_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3963__A2 _3960_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2799__A _2799_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2829_ _2829_/A _2846_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_351 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4496__RESET_B _2300_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_546 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4425__RESET_B _2385_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_139 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_419 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_590 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3423__A _3414_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_633 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4474__SET_B _2326_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_240 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_666 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_508 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_12 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3142__B _3151_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_390 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4254__A _3388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_533 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_577 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4404__D _4404_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3954__A2 _3952_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_82 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3706__A2 _3705_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2502__A _2497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3317__B _3316_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_110 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3333__A _3330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3890__A1 _4542_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2693__A2 _2691_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_636 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_124 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_349 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3052__B _3051_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_488 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_522 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_563 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_393 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4164__A _4585_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3801_ _3707_/A _2639_/X _3802_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_60_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_227 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_104 VGND VPWR sky130_fd_sc_hd__fill_2
X_3732_ _3726_/X _3669_/C _3719_/X _3731_/Y _3732_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_13_290 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_137 VGND VPWR sky130_fd_sc_hd__fill_1
X_3663_ _3508_/A _3437_/B _3663_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2412__A _2411_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3508__A _3508_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2614_ _4050_/A _4033_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_3594_ _2857_/A _3589_/X _3596_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3227__B _3375_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2545_ _2544_/X _2546_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4107__C1 _4106_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_387 VGND VPWR sky130_fd_sc_hd__decap_8
X_2476_ _2475_/X _2476_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_4215_ _4213_/Y _4215_/B _4216_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_95_260 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3243__A _2954_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2785__C _2785_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_614 VGND VPWR sky130_fd_sc_hd__decap_3
X_4146_ _4137_/B _4146_/B _4620_/D _4147_/C VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_28_305 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4452__CLK _4450_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_636 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_157 VGND VPWR sky130_fd_sc_hd__decap_4
X_4077_ utmi_data_out_o[4] _4076_/X _4079_/B VGND VPWR sky130_fd_sc_hd__nor2_4
X_3028_ _3015_/X _3016_/Y _3071_/A _3120_/B _3028_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_64_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_382 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_249 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_25 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2322__A _2318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3418__A _3427_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4606__RESET_B _2169_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_404 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3137__B _3207_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_227 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4249__A _4249_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4113__A2 _4111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3321__B1 _3319_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_603 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3153__A _3153_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_124 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_455 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2992__A _2944_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_488 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_511 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3600__B _3589_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_503 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_98 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_536 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2813__B1_N _2810_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3328__A _3563_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4325__CLK _4325_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2232__A _2236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4347__RESET_B _2478_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_170 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_264 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2589__D _2588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3047__B _3008_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2330_ _2330_/A _2330_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_216 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_205 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4475__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_346 VGND VPWR sky130_fd_sc_hd__decap_4
X_2261_ _2261_/A _2261_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4159__A _4143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3312__B1 _2986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3063__A _3010_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4000_ _3999_/Y _3994_/B _3962_/Y _3981_/X _4000_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_65_411 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_102 VGND VPWR sky130_fd_sc_hd__fill_2
X_2192_ _2188_/X _2192_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3700__A2_N _3699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_628 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2407__A _2408_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3510__B _3513_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_193 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4040__A1 _4562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3715_ _3713_/A _3715_/B _3715_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_107_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3238__A _2886_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3646_ _3528_/C _3528_/D _3498_/C _3528_/B _3646_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_115_630 VGND VPWR sky130_fd_sc_hd__fill_2
X_3577_ _3547_/A _3583_/B _3578_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_140 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_503 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2796__B _2796_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2528_ _2527_/Y _2525_/X _2528_/C _2528_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_102_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_547 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_15 VGND VPWR sky130_fd_sc_hd__decap_6
X_2459_ _2456_/A _2459_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_603 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3854__A1 _4527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4219__D _4219_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4129_ _2736_/X _4119_/X _4128_/X _4129_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_29_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_252 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_414 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_617 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2317__A _2324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_75 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_536 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3909__A2 _3897_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_193 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4348__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_569 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3148__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4498__CLK _4450_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_536 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_688 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4098__A1 _3955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_455 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3611__A outport_data_o[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_639 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3330__B _2860_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2872__D _2872_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_330 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2227__A _2228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4599__RESET_B _2177_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2820__A2 _2819_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_683 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4528__RESET_B _2262_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_366 VGND VPWR sky130_fd_sc_hd__fill_1
X_3500_ _3516_/B _3512_/B VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4161__B _4158_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3058__A _3359_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4480_ _3751_/X _3711_/B _2319_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_7_584 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_449 VGND VPWR sky130_fd_sc_hd__fill_2
X_3431_ _3498_/C _3556_/B _3431_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3208__D _3207_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3362_ _3397_/A _3358_/X _3362_/C _3362_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3505__B _3512_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2313_ _2314_/A _2313_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_143 VGND VPWR sky130_fd_sc_hd__fill_2
X_3293_ _3293_/A _3275_/B _3293_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3836__A1 utmi_rxvalid_i VGND VPWR sky130_fd_sc_hd__diode_2
X_2244_ _2241_/A _2244_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3224__C _3167_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_455 VGND VPWR sky130_fd_sc_hd__decap_3
X_2175_ _2177_/A _2175_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3521__A _2866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_200 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_458 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2811__A2 _2810_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_694 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4013__B2 _4012_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_16 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_254 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4502__D _3815_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4071__B _4072_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_265 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3772__B1 _3695_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_298 VGND VPWR sky130_fd_sc_hd__fill_2
X_3629_ _3612_/A _3627_/X _3628_/X _3629_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_88_300 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2600__A _2628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_666 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_230 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_444 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3431__A _3498_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_550 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_285 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4246__B _4235_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_127 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3150__B _3105_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_661 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_609 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_67 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_683 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4262__A _4610_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_642 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_199 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4412__D _4412_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_348 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3763__B1 _2659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3028__D _3120_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3606__A _3415_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2510__A _2159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2867__D _2866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_377 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_208 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4513__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_712 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3341__A _2857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3060__B _3038_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_553 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_90 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VPWR sky130_fd_sc_hd__decap_3
X_3980_ utmi_txready_i _3980_/B _3980_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2931_ _2930_/X _2972_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4243__B2 _4260_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4362__RESET_B _2459_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4172__A _4587_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2862_ _2862_/A _4405_/Q _4404_/Q _4407_/Q _2862_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_87_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_4601_ _4222_/X _4116_/D _2175_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_30_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_2793_ _2636_/A _2790_/X _2791_/Y _2792_/Y _2793_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XANTENNA__3754__B1 _3753_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4532_ _3866_/X _4532_/Q _2257_/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4322__D _4322_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_62 VGND VPWR sky130_fd_sc_hd__fill_2
X_4463_ _4525_/Q outport_data_o[5] _2340_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3516__A _3516_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2420__A _2419_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3414_ _3414_/A _3508_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_4394_ _3562_/Y _3559_/A _2421_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2777__D _2776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_141 VGND VPWR sky130_fd_sc_hd__fill_2
X_3345_ _3337_/Y _3344_/X _3345_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_112_496 VGND VPWR sky130_fd_sc_hd__fill_2
X_3276_ _3243_/B _2969_/X _3276_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3809__A1 _2641_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_509 VGND VPWR sky130_fd_sc_hd__fill_2
X_2227_ _2228_/A _2227_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3251__A _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_594 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_222 VGND VPWR sky130_fd_sc_hd__decap_4
X_2158_ _2252_/A _2159_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_296 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4066__B _4066_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_414 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_480 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_318 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3129__C _3119_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_268 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3426__A _3528_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2330__A _2330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_631 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_664 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3145__B _3144_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4536__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_697 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_185 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_369 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4257__A _4257_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3161__A _3161_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_296 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4407__D _4407_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4225__A1 _4224_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_447 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_469 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4225__B2 _4219_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_653 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2505__A _2504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_185 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_81 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_189 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3200__A2 _3014_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3336__A _2896_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2240__A _2241_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_362 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_100 VGND VPWR sky130_fd_sc_hd__fill_2
X_3130_ _3029_/X _3041_/X _3227_/D _3066_/A _3130_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__2894__B _2871_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_590 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3267__A2 _3265_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3071__A _3071_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4167__A _4197_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3061_ _3060_/X _3061_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_82_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_222 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_211 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4543__RESET_B _2243_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4317__D _2833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3221__D _3220_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_480 VGND VPWR sky130_fd_sc_hd__decap_8
X_3963_ _2605_/X _3960_/Y _3961_/X _2581_/X _3962_/Y _3963_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_3894_ _4544_/Q _3883_/X _3893_/X _4544_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__2415__A _2411_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2914_ _2914_/A _3241_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_269 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3975__B1 _2611_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_461 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4409__CLK _4410_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2845_ _4323_/Q _2829_/A _2844_/X _2845_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3727__B1 _3705_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4515_ _3829_/Y _3822_/A _2277_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_533 VGND VPWR sky130_fd_sc_hd__fill_2
X_2776_ _2771_/X _2772_/X _2776_/C _2775_/X _2776_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_105_717 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3246__A _3246_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2950__B2 _2949_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4446_ _4446_/D _4446_/Q _2359_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4559__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2150__A rst_i VGND VPWR sky130_fd_sc_hd__diode_2
X_4377_ _3655_/Y _3653_/A _2442_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3328_ _3563_/A _3329_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_358 VGND VPWR sky130_fd_sc_hd__decap_12
X_3259_ _3251_/X _3257_/X _3258_/X _4328_/Q _3248_/X _3260_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_85_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4077__A utmi_data_out_o[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_701 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_488 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_380 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3412__C _3411_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_553 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_406 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2325__A _2330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4434__SET_B _2373_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3718__B1 _3704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_627 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_656 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_137 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_409 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_66 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_472 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_314 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3603__B _3589_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_336 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3249__A2 _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_166 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_317 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_65 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_575 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_556 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2235__A _2236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4153__C _4147_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_409 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_258 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_421 VGND VPWR sky130_fd_sc_hd__fill_2
X_2630_ _2629_/X _2670_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_465 VGND VPWR sky130_fd_sc_hd__decap_4
X_2561_ _2560_/X _4278_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3066__A _3066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_225 VGND VPWR sky130_fd_sc_hd__decap_12
X_2492_ _2495_/A _2492_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4300_ _2526_/C _4299_/Y _2684_/X _4300_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_5_682 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4600__D _4221_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_258 VGND VPWR sky130_fd_sc_hd__fill_2
X_4231_ _2908_/C _3238_/C _4231_/C _2911_/B _4250_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_4_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_420 VGND VPWR sky130_fd_sc_hd__decap_3
X_4162_ _4187_/D _4158_/X _4163_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3513__B _3513_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_615 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_4093_ _3969_/Y _4016_/Y _4568_/Q utmi_data_out_o[6] _4093_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3113_ _3048_/Y _3098_/Y _3119_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_95_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_626 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_199 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_3044_ _3359_/B _3043_/X _3044_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_82_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_361 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_523 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_575 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_383 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_534 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_225 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3948__B1 _2611_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3946_ _2581_/A _3944_/X _3945_/X _2604_/X _4557_/Q _3946_/X VGND VPWR sky130_fd_sc_hd__o32a_4
X_3877_ _4545_/Q _3877_/B _3877_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3963__A3 _3961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2799__B _2796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4381__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2828_ _2557_/X _2910_/B _4316_/Q _2829_/A VGND VPWR sky130_fd_sc_hd__o21a_4
X_2759_ _4468_/Q _2548_/A _4469_/Q _2762_/C VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_3_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4510__D _4511_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_4429_ _3450_/Y _4429_/Q _2379_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4125__B1 _3980_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3704__A _3704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_431 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_252 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4465__RESET_B _2336_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_144 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_285 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_704 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_692 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2772__A1_N _4610_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4254__B _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_545 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_56 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_402 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3954__A3 _3953_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4270__A _4270_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3167__A1 _3205_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4420__D _4420_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3614__A outport_data_o[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_674 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_280 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2678__B1 _2654_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3333__B _3332_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3890__A2 _3883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_412 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_648 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_339 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_467 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_169 VGND VPWR sky130_fd_sc_hd__decap_12
X_3800_ _2601_/X _3785_/X _4496_/Q _2659_/X _3792_/A _4496_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_60_364 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_342 VGND VPWR sky130_fd_sc_hd__fill_2
X_3731_ _3724_/A _3729_/Y _3730_/X _3731_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_20_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_639 VGND VPWR sky130_fd_sc_hd__decap_12
X_3662_ _3662_/A _3430_/A _3661_/X _3662_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__4180__A _4180_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4480__SET_B _2319_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3593_ _3585_/X _3593_/B _3592_/X _3593_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_2613_ _2552_/X _2566_/X _2612_/X _4435_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__4330__D _4330_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2544_ _2534_/Y _2537_/X _2540_/X _2543_/X _2544_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3227__C _3011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_322 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4107__B1 _4033_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_377 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3524__A _2863_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2475_ _2496_/A _2475_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_228 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_431 VGND VPWR sky130_fd_sc_hd__fill_2
X_4214_ _2534_/Y _2714_/X _4213_/Y _4214_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_95_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3243__B _3243_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2785__D _4450_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_442 VGND VPWR sky130_fd_sc_hd__fill_2
X_4145_ _4146_/B _4137_/X _4147_/B VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_68_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_626 VGND VPWR sky130_fd_sc_hd__fill_2
X_4076_ _4011_/Y _4075_/X _4011_/Y _4075_/X _4076_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_106 VGND VPWR sky130_fd_sc_hd__fill_2
X_3027_ _4355_/Q _3120_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2841__B1 _2840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_16 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_545 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4505__D _3821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_567 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_578 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_217 VGND VPWR sky130_fd_sc_hd__decap_3
X_3929_ _4555_/Q _3929_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_109_127 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4090__A utmi_data_out_o[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_311 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3137__C _3136_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_333 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_438 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3434__A _2902_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_52 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3321__A1 _3234_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3153__B _3150_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_475 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_615 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2992__B _2985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_607 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4265__A _4265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_501 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4415__D _4415_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_386 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_93 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3609__A _3612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2513__A _2159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_609 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_193 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4387__RESET_B _2430_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2899__B1 _2898_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3047__C _3039_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_7 VGND VPWR sky130_fd_sc_hd__fill_1
X_2260_ _2253_/A _2261_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_239 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4316__RESET_B _2513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_358 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3312__B2 _3248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3312__A1 _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4159__B _4157_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_20 VGND VPWR sky130_fd_sc_hd__decap_12
X_2191_ _2188_/X _2191_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_92_231 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_467 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4175__A _4197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3076__B1 _3176_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_383 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4325__D _3323_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4040__A2 _4037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_559 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_414 VGND VPWR sky130_fd_sc_hd__fill_2
X_3714_ _3708_/X _3671_/X _3704_/X _3713_/X _4473_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3519__A _3547_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2423__A _2419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3238__B _2906_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_108 VGND VPWR sky130_fd_sc_hd__decap_12
X_3645_ _3662_/A _3643_/X _3644_/X _3645_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_20_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_3576_ _2855_/A _3566_/B _3576_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_2527_ _2522_/X _2527_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_114_185 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3254__A _2917_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_537 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2796__C _2793_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2458_ _2456_/A _2458_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2389_ _2396_/A _2391_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_581 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3854__A2 _3841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_242 VGND VPWR sky130_fd_sc_hd__fill_2
X_4128_ _2575_/C _4127_/X _3979_/X _4128_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_29_648 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4085__A _4079_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4059_ _4561_/Q _4058_/X _4059_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_71_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_43 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2814__B1 _2813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_353 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_548 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3429__A _3429_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2333__A _2337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3148__B _3143_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_257 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_174 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3164__A _3160_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4098__A2 _4039_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_710 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_380 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_294 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3611__B _3587_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2508__A _2504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_618 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3330__C _3329_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2805__B1 _2635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_695 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_301 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2243__A _2241_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2569__C1 _2705_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_389 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3230__B1 _2850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_530 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3058__B _3360_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4442__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3430_ _3430_/A _3556_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3361_ _2907_/X _3361_/B _3361_/C _3362_/C VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_112_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_100 VGND VPWR sky130_fd_sc_hd__fill_2
X_2312_ _2314_/A _2312_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4592__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_3292_ _3279_/A _3292_/B _3292_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3836__A2 _4519_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2243_ _2241_/A _2243_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_581 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3802__A _3802_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3224__D _3224_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_220 VGND VPWR sky130_fd_sc_hd__fill_2
X_2174_ _2166_/X _2177_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3521__B _3513_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2418__A _2419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_467 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_595 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_223 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2153__A _2155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_28 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3772__B2 _3771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3628_ outport_data_o[2] _3625_/B _3628_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_483 VGND VPWR sky130_fd_sc_hd__decap_4
X_3559_ _3559_/A _3566_/B _3562_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_103_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_47 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2328__A _2330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3431__B _3556_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_456 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4246__C _4239_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_139 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3150__C _3350_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_97 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_695 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4465__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_156 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_323 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_334 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_356 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3159__A _3148_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3776__A2_N _3771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3212__B1 _3412_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3763__B2 _2660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2998__A _2997_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3622__A outport_data_o[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_404 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2238__A _2238_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2970__A2_N _2969_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_297 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_286 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_437 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4015__A1_N _4011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_651 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3060__C _3039_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2930_ _2930_/A _2948_/A _2930_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_43_470 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_481 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_621 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_643 VGND VPWR sky130_fd_sc_hd__fill_2
X_2861_ _2860_/X _2861_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4603__D _4603_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4600_ _4221_/X _4116_/C _2176_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_30_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3069__A _3046_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_687 VGND VPWR sky130_fd_sc_hd__fill_2
X_2792_ _2804_/A _2691_/A _2636_/A _2792_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_698 VGND VPWR sky130_fd_sc_hd__decap_4
X_4531_ _3864_/X _4531_/Q _2258_/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3754__A1 _3745_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4331__RESET_B _2497_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4462_ _4524_/Q outport_data_o[4] _2341_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2701__A _2701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3516__B _3516_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3413_ _3413_/A _3657_/D _3414_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_98_632 VGND VPWR sky130_fd_sc_hd__fill_1
X_4393_ _4393_/D _4393_/Q _2422_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_97_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_507 VGND VPWR sky130_fd_sc_hd__fill_2
X_3344_ _3340_/X _3342_/X _3343_/Y _3344_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_100_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_315 VGND VPWR sky130_fd_sc_hd__decap_8
X_3275_ _2926_/A _3275_/B _3275_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3532__A _3503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3809__A2 _3803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4338__CLK _4430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2226_ _2228_/A _2226_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_231 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_510 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_2157_ _2155_/A _2157_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_81_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_543 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4488__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_492 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4419__RESET_B _2392_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4513__D utmi_rxactive_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_164 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_715 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3129__D _3181_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_214 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3707__A _3707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2611__A _2610_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_453 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_529 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_518 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3442__A _3424_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_540 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4257__B _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3681__B1 _3680_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_532 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_415 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_598 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4273__A _4368_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4225__A2 _4216_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_61 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_481 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4423__D _4423_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_676 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_113 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_658 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3617__A _3616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2521__A _4228_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_707 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3336__B _4375_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_217 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_291 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_197 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2894__C _2853_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3352__A _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3060_ _3007_/X _3038_/Y _3039_/Y _3009_/Y _3060_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3267__A3 _3266_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_679 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_551 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3071__B _4355_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4167__B _4167_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_418 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4583__RESET_B _2196_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3975__A1 _2572_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_492 VGND VPWR sky130_fd_sc_hd__decap_8
X_3962_ _4559_/Q _3962_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3893_ utmi_data_in_i[0] _3895_/B _3893_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4333__D _3284_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2913_ _3319_/A _2913_/B _2914_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3975__B2 _3974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4512__RESET_B _2280_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2844_ inport_data_i[6] _2846_/B _2844_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3727__A1 _3670_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3727__B2 _3702_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_545 VGND VPWR sky130_fd_sc_hd__decap_4
X_4514_ _3828_/X _4514_/Q _2278_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3527__A _3508_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2431__A _2431_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2775_ _4236_/A _2773_/Y _4266_/A _4494_/Q _2775_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_578 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_589 VGND VPWR sky130_fd_sc_hd__fill_2
X_4445_ _4308_/X _4445_/Q _2361_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4376_ _3652_/Y _4376_/Q _2443_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_98_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_451 VGND VPWR sky130_fd_sc_hd__decap_6
X_3327_ _3559_/A _3327_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3262__A _4329_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_434 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_3258_ _4328_/Q _3266_/B _3258_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_478 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_562 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4077__B _4076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4508__D _4508_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_329 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_510 VGND VPWR sky130_fd_sc_hd__decap_8
X_2209_ _2252_/A _2238_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_584 VGND VPWR sky130_fd_sc_hd__fill_2
X_3189_ _3068_/X _3144_/X _3189_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_26_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_351 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2606__A _2575_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_259 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3718__A1 _3708_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3437__A _3503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2341__A _2345_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4503__CLK _4450_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_283 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_101 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4268__A _4265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3172__A _3110_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_616 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3249__A3 _3247_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_307 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4418__D _3474_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_212 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3900__A utmi_data_in_i[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2516__A _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_568 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_484 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2955__A1_N _2954_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3347__A _3347_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2251__A _2248_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2560_ _2559_/X _2560_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2491_ _2495_/A _2491_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_672 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3066__B _3065_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_237 VGND VPWR sky130_fd_sc_hd__decap_6
X_4230_ _4247_/A _4276_/B _4605_/D VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_5_694 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_613 VGND VPWR sky130_fd_sc_hd__decap_12
X_4161_ _4187_/D _4158_/X _4161_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_4_64 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_112 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3082__A _4358_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4178__A _4186_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_156 VGND VPWR sky130_fd_sc_hd__fill_2
X_4092_ _3947_/A _4056_/X _4033_/A _4091_/Y _4092_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_3112_ _3112_/A _3112_/B _3190_/C _3111_/X _3112_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4328__D _4328_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3043_ _3031_/X _3105_/D _3015_/X _3043_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3810__A _3810_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_392 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4440__SET_B _2366_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_351 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2426__A _2431_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_237 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_clk_i clkbuf_3_7_0_clk_i/X clkbuf_5_30_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_51_568 VGND VPWR sky130_fd_sc_hd__fill_1
X_3945_ _4347_/Q _3417_/D _3945_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3948__B2 _4046_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3948__A1 _2571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4070__B1 _4012_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4526__CLK _4539_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_270 VGND VPWR sky130_fd_sc_hd__fill_2
X_3876_ _4536_/Q _3869_/X _3875_/X _3876_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_31_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_320 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3257__A _3265_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2827_ _4467_/Q _2796_/A _2783_/Y _2827_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__2161__A _2163_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2758_ _4050_/A _4443_/Q _2628_/C _4445_/Q _2762_/B VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_117_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_504 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_397 VGND VPWR sky130_fd_sc_hd__decap_8
X_2689_ _3713_/A _2689_/B _2689_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_4428_ _3446_/Y _4428_/Q _2380_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4125__A1 _2577_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_721 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_48 VGND VPWR sky130_fd_sc_hd__fill_2
X_4359_ _3373_/Y _4359_/Q _2463_/X _4334_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4088__A utmi_data_out_o[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_59 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_627 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_510 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3720__A _3720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_587 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2336__A _2337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_226 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_237 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_590 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_432 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4270__B _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_465 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_342 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3167__A2 _3088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_364 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_631 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3614__B _3587_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_292 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2678__A1 _2673_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2678__B2 _2677_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_432 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_443 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_605 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3630__A _3415_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_137 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_690 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_351 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4549__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2246__A _2248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_693 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_170 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_535 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4576__SET_B _2204_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_3730_ _3730_/A _3730_/B _3730_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_60_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_270 VGND VPWR sky130_fd_sc_hd__fill_2
X_3661_ _3528_/C _3498_/B _3661_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3592_ outport_data_o[0] _3592_/B _3592_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_70_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4611__D _4268_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_2612_ _2611_/X _2554_/X _2612_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2543_ _3808_/A _3806_/A _4502_/Q _4503_/Q _2543_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3805__A _3804_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3227__D _3227_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4107__A1 _3964_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3524__B _3513_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_2474_ _2472_/A _2474_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3866__B1 _3865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_4213_ _2711_/X _4213_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_68_465 VGND VPWR sky130_fd_sc_hd__decap_4
X_4144_ _4144_/A _4146_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_329 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3540__A _4405_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4075_ _3941_/Y _4565_/Q _3941_/Y _4565_/Q _4075_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_479 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_619 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4291__B1 _4288_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_351 VGND VPWR sky130_fd_sc_hd__decap_4
X_3026_ _3021_/X _3105_/D _3350_/C _3359_/B _3026_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_51_321 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2841__A1 _4321_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2156__A _2155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_365 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_557 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_387 VGND VPWR sky130_fd_sc_hd__fill_2
X_3928_ _3928_/A _2560_/X _3928_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_590 VGND VPWR sky130_fd_sc_hd__decap_8
X_3859_ _4537_/Q _3859_/B _3859_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_109_106 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4090__B _4090_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4521__D _3840_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3715__A _3713_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3857__B1 _3856_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3434__B _3434_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_432 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3321__A2 _2992_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3153__C _3151_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_35 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_13 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_638 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4615__RESET_B _2156_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_595 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3450__A _3424_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2992__C _2988_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4265__B _4263_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_107 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_630 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_395 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_398 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4281__A _4281_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_61 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3609__B _3607_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_723 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4431__D _3458_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3625__A outport_data_o[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2899__A1 _2891_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_288 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3047__D _3010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_505 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3848__B1 _3847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3312__A2 _3310_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2190_ _2188_/X _2190_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4159__C _4158_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_262 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4356__RESET_B _2466_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4371__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_148 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3360__A _3360_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_254 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_619 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4175__B _4178_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3076__A1 _3036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4606__D _4247_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_343 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_685 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4025__B1 _4024_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_404 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_590 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4191__A _4185_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2704__A _2704_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3713_ _3713_/A _3713_/B _3713_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3519__B _3516_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2587__B1 _4342_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_448 VGND VPWR sky130_fd_sc_hd__fill_2
X_3644_ outport_data_o[7] _3617_/X _3644_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4341__D _3317_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3238__C _3238_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3535__A _3506_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3575_ _3581_/A _3573_/Y _3574_/X _3575_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_115_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_654 VGND VPWR sky130_fd_sc_hd__fill_2
X_2526_ _2522_/X _2525_/X _2526_/C _2531_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_102_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3254__B _3266_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2796__D _2795_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2771__A1_N _4266_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2457_ _2456_/A _2457_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_197 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_348 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_28 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_39 VGND VPWR sky130_fd_sc_hd__fill_2
X_2388_ _2388_/A _2388_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_571 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_616 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3270__A _4331_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_370 VGND VPWR sky130_fd_sc_hd__fill_1
X_4127_ _2612_/X _4127_/B _4127_/C _4126_/X _4127_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__4085__B _4083_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4058_ _3918_/Y utmi_data_out_o[1] _3918_/Y _3925_/X _4058_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4516__D _3831_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2814__A1 _2803_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3009_ _4359_/Q _3009_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_674 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_140 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_376 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_48 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_509 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2614__A _4050_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3775__C1 _3774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3148__C _3108_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_571 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3445__A _3510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_665 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_52 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3164__B _3163_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_668 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4394__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_582 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_273 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_413 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4276__A _2516_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3180__A _3136_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_660 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4426__D _4426_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_671 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2805__A1 _2785_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_343 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_482 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2524__A _2522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3230__A1 _3229_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2569__B1 _2566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_542 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3058__C _3021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_564 VGND VPWR sky130_fd_sc_hd__fill_2
X_3360_ _3360_/A _3360_/B _3361_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4537__RESET_B _2250_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_613 VGND VPWR sky130_fd_sc_hd__decap_3
X_2311_ _2314_/A _2311_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_668 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_335 VGND VPWR sky130_fd_sc_hd__fill_2
X_3291_ _3280_/X _3289_/X _3290_/X _3289_/A _3277_/X _3292_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
X_2242_ _2241_/A _2242_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_530 VGND VPWR sky130_fd_sc_hd__fill_2
X_2173_ _2168_/A _2173_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4186__A _4164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_660 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_287 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4336__D _3296_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2434__A _2434_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_346 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3265__A _3265_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3627_ _2880_/A _3620_/B _3627_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2980__B1 _2979_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3558_ _3583_/B _3566_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_602 VGND VPWR sky130_fd_sc_hd__fill_2
X_2509_ _2504_/A _2509_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_103_646 VGND VPWR sky130_fd_sc_hd__fill_2
X_3489_ _3547_/A _3486_/B _3490_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_76_508 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_571 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_468 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_202 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_276 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4246__D _4245_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_438 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_427 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_65 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3150__D _3150_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_279 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_124 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_471 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2344__A _2345_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_157 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3159__B _3153_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3212__A1 _3210_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_390 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_40 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_62 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3175__A _3153_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2723__B1 _2602_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3622__B _3625_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2519__A _2518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_533 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_70 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3060__D _3009_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_674 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2254__A _2258_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2860_ _2855_/X _2857_/X _2860_/C _2860_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_70_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_132 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3069__B _3038_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2791_ _2691_/B _2791_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_716 VGND VPWR sky130_fd_sc_hd__decap_8
X_4530_ _4530_/D _4530_/Q _2259_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3754__A2 _3752_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_215 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2962__B1 _2961_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4461_ _4523_/Q outport_data_o[3] _2342_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2701__B _2700_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_383 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_75 VGND VPWR sky130_fd_sc_hd__fill_2
X_3412_ _3412_/A _3412_/B _3411_/Y _3412_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3085__A _3085_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4371__RESET_B _2449_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4392_ _4392_/D _4392_/Q _2423_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3343_ _3330_/X _3340_/X _3332_/X _3343_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3274_ _3246_/A _3275_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3532__B _3541_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_338 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2429__A _2431_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_722 VGND VPWR sky130_fd_sc_hd__decap_3
X_2225_ _2228_/A _2225_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_54_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_2156_ _2155_/A _2156_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_449 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2164__A _2163_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_17 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_21_0_clk_i_A clkbuf_5_21_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_622 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_633 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_143 VGND VPWR sky130_fd_sc_hd__fill_2
X_2989_ _3314_/A _2986_/Y _2989_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_176 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2953__B1 _2900_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4459__RESET_B _2344_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_515 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3723__A _3670_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_465 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_498 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3442__B _3439_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2339__A _2339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_530 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3130__B1 _3227_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3681__B2 _4474_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_371 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4432__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_585 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_235 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_577 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4273__B _4263_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4225__A3 _4214_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_633 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_441 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_430 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4582__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_132 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_474 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2802__A _2626_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3197__B1 _3114_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2944__B1 _3455_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_719 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3336__C _3335_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_353 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3914__A1_N _2571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3633__A _3662_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_143 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_284 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2249__A _2248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_135 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2894__D _2878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_338 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3071__C _3023_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4167__C _4166_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_279 VGND VPWR sky130_fd_sc_hd__fill_1
X_3961_ _3216_/A _4278_/C _3961_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2912_ _2912_/A _2913_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4614__D _4614_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3892_ _4543_/Q _3883_/X _3891_/X _3892_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_92_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_290 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3975__A2 _3973_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_452 VGND VPWR sky130_fd_sc_hd__decap_6
X_2843_ _4322_/Q _2831_/X _2842_/X _4322_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3727__A2 _3679_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2774_ _4608_/Q _2766_/Y _4236_/A _2773_/Y _2776_/C VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3808__A _3808_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2712__A _4353_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_513 VGND VPWR sky130_fd_sc_hd__decap_12
X_4513_ utmi_rxactive_i _4513_/Q _2279_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_681 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4552__RESET_B _2233_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_229 VGND VPWR sky130_fd_sc_hd__decap_8
X_4444_ _2742_/Y _4228_/B _2362_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3130__A2_N _3041_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4375_ _3649_/Y _4375_/Q _2444_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3543__A _3543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_463 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_11_0_clk_i clkbuf_3_5_0_clk_i/X clkbuf_5_22_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_3326_ _3347_/A _3325_/X _3347_/A _3325_/X _3326_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3262__B _3266_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_496 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_485 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4455__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_327 VGND VPWR sky130_fd_sc_hd__decap_4
X_3257_ _3265_/A _3257_/B _3257_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2159__A _2159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_596 VGND VPWR sky130_fd_sc_hd__decap_12
X_3188_ _3188_/A _3220_/C _3188_/C _3188_/D _3191_/C VGND VPWR sky130_fd_sc_hd__or4_4
X_2208_ _2206_/A _2208_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_94_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4076__A1_N _4011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4524__D _3848_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_396 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_216 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2606__B _4437_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_636 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_463 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3718__A2 _3683_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_607 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3179__B1 _3178_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3437__B _3437_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_117 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4014__A1_N utmi_data_out_o[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3728__A2_N _3727_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_441 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_312 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3453__A _3516_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3351__B1 _3360_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_367 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2984__A2_N _3303_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4268__B _4266_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3172__B _3018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_56 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_680 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_714 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3900__B _3904_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_224 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_341 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_717 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_268 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_205 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4434__D _2617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4328__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3628__A outport_data_o[2] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2532__A _4489_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3347__B _3347_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_489 VGND VPWR sky130_fd_sc_hd__fill_2
X_2490_ _2495_/A _2490_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_662 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4478__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_194 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_400 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3363__A _3363_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4160_ _4160_/A _4187_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_122_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_433 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_625 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4609__D _4609_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3082__B _4359_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4178__B _4178_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3111_ _3150_/D _3107_/Y _3108_/X _3110_/Y _3111_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_4091_ _4079_/A _4091_/B _4090_/X _4091_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_95_477 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_680 VGND VPWR sky130_fd_sc_hd__fill_2
X_3042_ _3041_/X _3219_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3810__B _3805_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_544 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4194__A _4591_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2707__A _2707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_514 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_503 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_205 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_683 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4344__D _4344_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3944_ _4321_/Q _3944_/B _3944_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3948__A2 _3946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_249 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4070__B2 _4069_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3875_ _4544_/Q _3877_/B _3875_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3538__A _3510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2442__A _2443_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2826_ _2825_/X _2826_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3257__B _3257_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_332 VGND VPWR sky130_fd_sc_hd__fill_2
X_2757_ _2716_/Y _2761_/A _2757_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2688_ _2673_/X _2674_/Y _2642_/X _2652_/X _2689_/B VGND VPWR sky130_fd_sc_hd__or4_4
X_4427_ _4427_/D _4427_/Q _2383_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4125__A2 _4124_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3273__A _3240_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_603 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_16 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_647 VGND VPWR sky130_fd_sc_hd__fill_2
X_4358_ _3368_/Y _4358_/Q _2464_/X _4334_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4088__B _4087_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4519__D _4519_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_658 VGND VPWR sky130_fd_sc_hd__fill_2
X_3309_ _3317_/A _3308_/Y _4339_/D VGND VPWR sky130_fd_sc_hd__nor2_4
X_4289_ _4497_/Q _4286_/X _2533_/X _4289_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_100_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_160 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_193 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_36 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4403__RESET_B _2411_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3448__A outport_data_o[3] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2352__A _2352_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_52 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_23 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4620__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_78 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4279__A _4277_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_621 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_593 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2678__A2 _2674_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_175 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4429__D _3450_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_71 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_511 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3911__A _3005_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_672 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2527__A _2522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_385 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2262__A _2261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_591 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_231 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_129 VGND VPWR sky130_fd_sc_hd__decap_8
X_3660_ _3660_/A _3498_/B _3660_/C _3660_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_9_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_275 VGND VPWR sky130_fd_sc_hd__fill_2
X_3591_ _3587_/X _3592_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_2611_ _2610_/Y _2611_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2542_ _4498_/Q _3806_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4107__A2 _4039_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2473_ _2472_/A _2473_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4189__A _4182_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4212_ _4210_/X _4211_/X _4212_/C _4212_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3093__A _3068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3866__A1 _4532_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_422 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_530 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4339__D _4339_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4143_ _4140_/Y _4143_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_83_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_639 VGND VPWR sky130_fd_sc_hd__fill_2
X_4074_ _4570_/Q _4056_/X _4050_/X _4073_/Y _4570_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3540__B _3543_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_138 VGND VPWR sky130_fd_sc_hd__fill_2
X_3025_ _3016_/Y _3359_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_71_609 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2437__A _2434_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_190 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4291__B2 _4290_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4291__A1 _2548_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3115__A1_N _3061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2841__A2 _2831_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_344 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3268__A _3268_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3927_ _4319_/Q _2585_/A _3927_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_3858_ _3824_/X _3859_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_17 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2172__A _2168_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2809_ _4514_/Q _2784_/A _2808_/X _2809_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_3789_ _3685_/X _3782_/X _3790_/B _4489_/Q _3786_/Y _4489_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_105_302 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2900__A _2900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3715__B _3715_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_37 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4099__A _4009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_8 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_327 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3857__A1 _3837_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_411 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_390 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3153__D _3153_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3731__A _3724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_628 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3450__B _3450_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2992__D _2991_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_127 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4265__C _4265_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2347__A _2352_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_653 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_569 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_366 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_73 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3178__A _3058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3609__C _3608_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3793__B1 _4527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3906__A utmi_data_in_i[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2810__A _2636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3625__B _3625_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2899__A2 _2892_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_208 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3848__A1 _4524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_539 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_338 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3312__A3 _3311_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4516__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3641__A outport_data_o[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3360__B _3360_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2257__A _2258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_609 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4175__C _4175_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3076__A2 _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4396__RESET_B _2419_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_620 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4325__RESET_B _2504_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_697 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4025__A1 _4022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2587__A1 _4316_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4191__B _4192_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3088__A _3087_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3712_ _3708_/X _4472_/Q _3704_/X _3711_/X _4472_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__2587__B2 _3417_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3643_ _3643_/A _3640_/B _3643_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3238__D _2907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_600 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3816__A _3816_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2720__A _2715_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3535__B _3541_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3574_ _3516_/A _3583_/B _3574_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_114_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_143 VGND VPWR sky130_fd_sc_hd__decap_4
X_2525_ _4487_/Q _2525_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2456_ _2456_/A _2456_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3551__A _3522_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2387_ _2388_/A _2387_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_241 VGND VPWR sky130_fd_sc_hd__decap_12
X_4126_ _4123_/X _4125_/X _2569_/X _4126_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_28_105 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3270__B _3266_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_233 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3684__A1_N _2660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_266 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2768__A2_N _4490_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2167__A _2166_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4057_ _3974_/Y _4017_/Y _3974_/A utmi_data_out_o[0] _4061_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4085__C _4085_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_108 VGND VPWR sky130_fd_sc_hd__fill_2
X_3008_ _4360_/Q _3008_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_37_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2814__A2 _2812_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_642 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_152 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4532__D _3866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3775__B1 _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3726__A _3708_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2630__A _2629_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3148__D _3228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3445__B _3437_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_677 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_636 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_625 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4539__CLK _4539_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_165 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3461__A outport_data_o[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_285 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_436 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4276__B _4276_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_116 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3180__B _3176_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_417 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2805__A2 _2804_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_50 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_322 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_94 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_377 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_494 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2524__B _2523_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4442__D _2550_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2569__A1 _2568_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_369 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3230__A2 _2916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_510 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3636__A _3662_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3058__D _3347_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2540__A _2532_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_2310_ _2324_/A _2314_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_3290_ _3243_/B _2976_/X _3290_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2241_ _2241_/A _2241_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_78_550 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3371__A _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_425 VGND VPWR sky130_fd_sc_hd__decap_12
X_2172_ _2168_/A _2172_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4577__RESET_B _2203_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4186__B _4186_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4506__RESET_B _2287_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4617__D _4296_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_299 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2715__A _2711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_336 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3757__B1 _3667_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4352__D _2996_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_358 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3546__A _4407_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2980__A1 _3297_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2450__A _2449_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3626_ _3612_/A _3626_/B _3625_/X _4379_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_115_452 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3265__B _3265_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3557_ _3557_/A _3583_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_2508_ _2504_/A _2508_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_658 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_124 VGND VPWR sky130_fd_sc_hd__fill_2
X_3488_ _3488_/A _3478_/B _3488_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3281__A _2928_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_550 VGND VPWR sky130_fd_sc_hd__fill_2
X_2439_ _2425_/A _2443_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4527__D _3854_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_255 VGND VPWR sky130_fd_sc_hd__fill_2
X_4109_ _4009_/X _4108_/B _4108_/X _4109_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_84_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_119 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_480 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_631 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2625__A _4449_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_48 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3159__C _3158_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3212__A2 _2999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3456__A outport_data_o[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_380 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4361__CLK _4334_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_524 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2360__A _2339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3175__B _3165_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2723__A1 _2707_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_433 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_336 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4287__A _2716_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3191__A _3136_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_542 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_704 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_233 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4437__D _2603_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_277 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_480 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2535__A _4504_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_461 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_280 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_111 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3069__C _3011_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2790_ _2694_/A _2790_/B _2790_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3366__A _3366_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_351 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_54 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2962__A1 _4329_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2270__A _2272_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4460_ _4522_/Q outport_data_o[2] _2343_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_362 VGND VPWR sky130_fd_sc_hd__decap_4
X_4391_ _3609_/X _3607_/A _2426_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3411_ _4392_/Q _3398_/B _3411_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_7_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3085__B _3085_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3342_ _2867_/A _3342_/B _3342_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_3273_ _3240_/A _3279_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4197__A _4197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_211 VGND VPWR sky130_fd_sc_hd__decap_3
X_2224_ _2238_/A _2228_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4340__RESET_B _2486_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2155_ _2155_/A _2155_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_255 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4347__D _3203_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_523 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2445__A _2443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_450 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4384__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_2988_ _3460_/A _2987_/X _3460_/A _2987_/X _2988_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__3276__A _3243_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_25_0_clk_i_A clkbuf_5_25_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_227 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2953__B2 _3265_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2180__A _2177_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3609_ _3612_/A _3607_/X _3608_/X _3609_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_89_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_601 VGND VPWR sky130_fd_sc_hd__decap_8
X_4589_ _4184_/Y _4182_/A _2189_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4499__RESET_B _2297_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3723__B _3723_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_99 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4428__RESET_B _2380_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3442__C _3441_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_520 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_211 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3130__B2 _3066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_361 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_299 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2355__A _2358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4244__A1_N _4610_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_111 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_605 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_689 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3197__A1 _3045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2802__B _2638_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3186__A _3186_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2944__B2 _2943_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_306 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3633__B _3633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_296 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3771__B1_N _3770_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_597 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3071__D _4357_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2265__A _2261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_589 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_567 VGND VPWR sky130_fd_sc_hd__fill_2
X_3960_ _4323_/Q _3960_/B _3960_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_90_386 VGND VPWR sky130_fd_sc_hd__decap_6
X_2911_ _4342_/Q _2911_/B _2912_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_3891_ _3891_/A _3895_/B _3891_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2842_ inport_data_i[5] _2846_/B _2842_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_486 VGND VPWR sky130_fd_sc_hd__fill_2
X_2773_ _4492_/Q _2773_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3808__B _3805_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2712__B _3417_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_525 VGND VPWR sky130_fd_sc_hd__decap_8
X_4512_ _4513_/Q _4512_/Q _2280_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_569 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_693 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3824__A _3824_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4443_ _2756_/X _4443_/Q _2363_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_98_431 VGND VPWR sky130_fd_sc_hd__fill_2
X_4374_ _4374_/D _3244_/B _2445_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4592__RESET_B _2185_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3543__B _3543_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4521__RESET_B _2270_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_615 VGND VPWR sky130_fd_sc_hd__decap_4
X_3325_ _3324_/X _3325_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_3256_ _3268_/A _3256_/B _4327_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_85_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_531 VGND VPWR sky130_fd_sc_hd__decap_12
X_2207_ _2206_/A _2207_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3187_ _3045_/X _3085_/B _3188_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_26_203 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_534 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_589 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_556 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2995__B1_N _2994_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2175__A _2177_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2606__C _2606_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4058__A2_N utmi_data_out_o[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2903__A _3455_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_615 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3179__A1 _3013_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4540__D _4540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_525 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_503 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4128__B1 _3979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4609__RESET_B _2164_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_76 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_58 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_36 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_252 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3453__B _3462_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3351__A1 _3359_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_125 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4268__C _4267_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_670 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4300__B1 _2684_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_394 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_383 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_534 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_364 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_375 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_83 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3628__B _3625_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2532__B _4488_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_497 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4450__D _4450_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_9 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3347__C _3325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3644__A outport_data_o[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_580 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3363__B _3325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_583 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_80 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3082__C _3007_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3110_ _3011_/X _3369_/A _3110_/C _3382_/A _3110_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_4_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_456 VGND VPWR sky130_fd_sc_hd__fill_2
X_4090_ utmi_data_out_o[6] _4090_/B _4090_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_95_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VPWR sky130_fd_sc_hd__fill_2
X_3041_ _3040_/X _3041_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_63_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2707__B _2706_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4055__C1 _4054_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_194 VGND VPWR sky130_fd_sc_hd__fill_1
X_3943_ _3943_/A utmi_data_out_o[3] VGND VPWR sky130_fd_sc_hd__buf_1
X_3874_ _4535_/Q _3869_/X _3873_/X _3874_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_31_261 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3538__B _3541_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2825_ _2620_/B _2800_/X _2825_/C _2824_/X _2825_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__4360__D _4360_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2756_ _2743_/X _2755_/X _2602_/X _2756_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_117_355 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3554__A _3554_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4422__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2687_ _3704_/A _2687_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4426_ _4426_/D _2902_/D _2384_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_200 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_423 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_28 VGND VPWR sky130_fd_sc_hd__decap_3
X_4357_ _3362_/Y _4357_/Q _2465_/X _4356_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4572__CLK _4574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_594 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_147 VGND VPWR sky130_fd_sc_hd__fill_2
X_3308_ _3251_/A _3306_/X _3307_/X _3306_/A _3248_/A _3308_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_4288_ _2760_/X _4287_/X _2533_/X _4288_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_73_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_169 VGND VPWR sky130_fd_sc_hd__fill_2
X_3239_ _3397_/A _3236_/X _3238_/X _3239_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_67_681 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4535__D _3874_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_49 VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_9_0_clk_i clkbuf_4_9_0_clk_i/A clkbuf_4_9_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_15_707 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_578 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_66 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3729__A _3730_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2633__A _4514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_581 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_412 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4443__RESET_B _2363_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3464__A _3464_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4279__B _4278_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_132 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2678__A3 _2661_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_136 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_670 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3911__B _2560_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_448 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2835__B1 _2834_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4445__D _4308_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_194 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3639__A _3662_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_389 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2543__A _3808_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_261 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4445__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_108 VGND VPWR sky130_fd_sc_hd__decap_4
X_3590_ _2867_/A _3589_/X _3593_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_2610_ _2610_/A _2610_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2541_ _4499_/Q _3808_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3374__A _3353_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2472_ _2472_/A _2472_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4595__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_509 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4189__B _4186_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4075__A1_N _3941_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4211_ _3987_/A _2704_/A _4211_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3866__A2 _3855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_542 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_456 VGND VPWR sky130_fd_sc_hd__fill_2
X_4142_ _4135_/X _4137_/X _4197_/A _4142_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_95_264 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_670 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2718__A _2716_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4073_ _4073_/A _4071_/Y _4072_/X _4073_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_28_309 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_448 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_681 VGND VPWR sky130_fd_sc_hd__fill_2
X_3024_ _3023_/Y _3350_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_64_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4291__A2 _2761_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4355__D _3349_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_673 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_386 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_364 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4013__A1_N utmi_data_out_o[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3549__A _3508_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2453__A _2425_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_3926_ _2552_/A _3918_/Y _3925_/X utmi_data_out_o[1] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3268__B _3268_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_721 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_581 VGND VPWR sky130_fd_sc_hd__decap_3
X_3857_ _3837_/A _3855_/X _3856_/X _3857_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_118_642 VGND VPWR sky130_fd_sc_hd__decap_4
X_2808_ _2636_/A _2803_/X _2807_/Y _2808_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_3788_ _2657_/X _3782_/X _3790_/B _4488_/Q _3786_/Y _3788_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_117_141 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2900__B _4420_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2739_ _2727_/X _2741_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_163 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3284__A _3279_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_419 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_358 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4099__B _4099_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4409_ _4409_/D _2865_/B _2404_/X _4410_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3857__A2 _3855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_33 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_542 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3731__B _3729_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2628__A _2694_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_607 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3450__C _3449_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4318__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_640 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_342 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_504 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_515 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_526 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_183 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4468__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3459__A _3660_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_378 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2363__A _2362_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_518 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3793__A1 _2522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3178__B _3047_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3793__B2 _3792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_253 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_620 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_653 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3906__B _3904_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2810__B _2810_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_62 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3194__A _2850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3848__A2 _3841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_485 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3641__B _3617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_415 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2538__A _4501_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_34 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_245 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2808__B1 _2807_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_470 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_312 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2273__A _2272_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3369__A _3369_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_356 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4025__A2 _4024_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_581 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3711_ _3713_/A _3711_/B _3711_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4365__RESET_B _2456_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2587__A2 _3960_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_439 VGND VPWR sky130_fd_sc_hd__fill_2
X_3642_ _3662_/A _3642_/B _3641_/X _3642_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3816__B _3805_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_634 VGND VPWR sky130_fd_sc_hd__decap_12
X_3573_ _2855_/B _3566_/B _3573_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2720__B _4278_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_667 VGND VPWR sky130_fd_sc_hd__decap_4
X_2524_ _2522_/X _2523_/Y _2524_/C _2524_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_88_529 VGND VPWR sky130_fd_sc_hd__decap_8
X_2455_ _2456_/A _2455_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3832__A _4518_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_540 VGND VPWR sky130_fd_sc_hd__decap_12
X_2386_ _2388_/A _2386_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3551__B _3544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_253 VGND VPWR sky130_fd_sc_hd__decap_12
X_4125_ _2577_/Y _4124_/X _3980_/B _4125_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_84_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2448__A _2449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_128 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_4056_ _4079_/A _4056_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_71_418 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4610__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3007_ _4361_/Q _3007_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_101_13 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_492 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_120 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3279__A _3279_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2183__A _2183_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_389 VGND VPWR sky130_fd_sc_hd__decap_4
X_3909_ _3891_/A _3897_/X _3908_/X _3909_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3775__A1 _3724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2911__A _4342_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_648 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_114 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_540 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_169 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_404 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2358__A _2358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_201 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4276__C _4275_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_234 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3180__C _3077_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_429 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_470 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_684 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_clk_i clkbuf_3_7_0_clk_i/A clkbuf_3_6_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_43_654 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_621 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_367 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3189__A _3068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_304 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2524__C _2524_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2569__A2 _2562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2821__A _2821_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_562 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3917__A _3916_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3636__B _3634_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_472 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_461 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2540__B _2539_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_599 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_315 VGND VPWR sky130_fd_sc_hd__decap_12
X_2240_ _2241_/A _2240_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_348 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3652__A _3581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3371__B _3342_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2268__A _2272_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_510 VGND VPWR sky130_fd_sc_hd__decap_8
X_2171_ _2168_/A _2171_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_610 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_481 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4546__RESET_B _2240_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2715__B _2714_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_153 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3099__A _3084_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3757__B2 _3668_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_214 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3827__A _3883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2731__A _2537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3546__B _3543_/B VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_8_0_clk_i clkbuf_5_9_0_clk_i/A _4509_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__2953__A1_N _2900_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3625_ outport_data_o[1] _3625_/B _3625_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2980__A2 _2935_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_420 VGND VPWR sky130_fd_sc_hd__decap_3
X_3556_ _3528_/A _3556_/B _3557_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_103_626 VGND VPWR sky130_fd_sc_hd__decap_4
X_2507_ _2504_/A _2507_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3487_ _3504_/A _3485_/Y _3486_/X _4422_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3562__A _3555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_158 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3281__B _3275_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2438_ _2434_/A _2438_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_702 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3693__B1 _2650_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_2369_ _2367_/X _2369_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2178__A _2177_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_404 VGND VPWR sky130_fd_sc_hd__decap_12
X_4108_ _4009_/X _4108_/B _4108_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2906__A _2899_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4039_ _3923_/Y _4039_/B _4039_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_112_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4543__D _3892_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_613 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_304 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_687 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_159 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3159__D _3119_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3737__A _3724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2641__A _4521_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4506__CLK _4450_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_503 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_442 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3175__C _3167_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2723__A2 _2722_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3472__A _3486_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4287__B _4286_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3191__B _3176_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3684__B1 _2660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_510 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_191 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_392 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_716 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2816__A _2815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_492 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_440 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_602 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4453__D _2631_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_60 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3069__D _3010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3647__A _4375_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_93 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_11 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2551__A _3925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3366__B _3343_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2962__A2 _2920_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4390_ _3605_/X _2858_/B _2427_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2767__A2_N _2765_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3410_ _4368_/Q _3394_/B _3412_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_98_624 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_613 VGND VPWR sky130_fd_sc_hd__fill_2
X_3341_ _2857_/A _3342_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_434 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_635 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_112 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3382__A _3382_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3272_ _3268_/A _3271_/Y _4331_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_97_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4197__B _4197_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_2223_ _2217_/X _2223_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_543 VGND VPWR sky130_fd_sc_hd__decap_4
X_2154_ _2155_/A _2154_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_93_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_587 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_267 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2726__A _3417_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_579 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4380__RESET_B _2438_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4529__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4363__D _3393_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_668 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3557__A _3557_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2987_ _2986_/A _2986_/B _2986_/Y _2987_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_21_156 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2461__A _2460_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3276__B _2969_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3608_ outport_data_o[5] _3592_/B _3608_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_401 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_9 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_29_0_clk_i_A clkbuf_5_29_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4588_ _4181_/Y _4176_/A _2190_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3539_ _3545_/A _3537_/Y _3539_/C _4404_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_107_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_635 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3292__A _3279_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_668 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4538__D _4538_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_554 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4468__RESET_B _2333_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_502 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_418 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2636__A _2636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_248 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_53 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4226__A2_N _4225_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_101 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_473 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3467__A _3483_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_189 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2371__A _2367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3197__A2 _3196_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3186__B _3216_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_366 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_123 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3633__C _3632_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4448__D _4448_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_583 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_159 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_340 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2546__A _2724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4082__B1 _4018_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_451 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_207 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_270 VGND VPWR sky130_fd_sc_hd__fill_2
X_2910_ _2560_/X _2910_/B _2911_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_3890_ _4542_/Q _3883_/X _3889_/X _3890_/X VGND VPWR sky130_fd_sc_hd__a21o_4
Xclkbuf_2_3_0_clk_i clkbuf_2_3_0_clk_i/A clkbuf_3_7_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_2841_ _4321_/Q _2831_/X _2840_/X _2841_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_31_465 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2281__A _2253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_2772_ _4610_/Q _2770_/Y _4612_/Q _2765_/Y _2772_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_498 VGND VPWR sky130_fd_sc_hd__decap_8
X_4511_ _4512_/Q _4511_/Q _2282_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_537 VGND VPWR sky130_fd_sc_hd__fill_2
X_4442_ _2550_/Y _2548_/A _2364_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_171 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3824__B utmi_rxvalid_i VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3896__B1 _3895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_410 VGND VPWR sky130_fd_sc_hd__decap_4
X_4373_ _3422_/X _2849_/A _2447_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3324_ _2913_/B _3322_/X _3324_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4001__A _2736_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3255_ _3251_/X _3253_/X _3254_/X _2917_/A _3248_/X _3256_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XANTENNA__4358__D _3368_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_510 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_448 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_543 VGND VPWR sky130_fd_sc_hd__fill_2
X_2206_ _2206_/A _2206_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3186_ _3186_/A _3216_/B _3186_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_66_384 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2456__A _2456_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4351__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_410 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2903__B _3460_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2191__A _2188_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3179__A2 _3177_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_559 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4128__A1 _2575_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_44 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_5_0_clk_i clkbuf_4_5_0_clk_i/A clkbuf_4_5_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_78_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_231 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3351__A2 _3347_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_498 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_627 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4565__SET_B _2218_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_297 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3750__A _3708_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4300__A1 _2526_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2366__A _2362_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_85 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4064__B1 _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3811__B1 _3810_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_432 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_270 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_454 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_476 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_95 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_295 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2532__C _2531_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_469 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3925__A _3925_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4103__A2_N _4102_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3878__B1 _3877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3644__B _3617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_697 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_686 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_540 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3082__D _3008_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3660__A _3660_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4374__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4319__RESET_B _2510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_619 VGND VPWR sky130_fd_sc_hd__fill_1
X_3040_ _4361_/Q _3038_/Y _3039_/Y _4359_/Q _3040_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2276__A _2277_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_310 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_696 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_376 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_527 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4055__B1 _4050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_229 VGND VPWR sky130_fd_sc_hd__fill_2
X_3942_ _2578_/X _3940_/X _2552_/X _3941_/Y _3943_/A VGND VPWR sky130_fd_sc_hd__o22a_4
X_3873_ _4543_/Q _3877_/B _3873_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2824_ _2821_/A _2788_/A _2796_/B _2823_/Y _2824_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_117_301 VGND VPWR sky130_fd_sc_hd__decap_4
X_2755_ _2715_/X _2745_/Y _2754_/Y _2755_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_117_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_2686_ _2684_/X _3713_/A _2785_/C _2666_/X _2670_/B _4450_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__3554__B _3544_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4425_ _4425_/D _3494_/A _2385_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4243__A1_N _4242_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4356_ _3357_/Y _4356_/Q _2466_/X _4356_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3307_ _3253_/A _2943_/X _3307_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3570__A _3513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_446 VGND VPWR sky130_fd_sc_hd__decap_12
X_4287_ _2716_/Y _4286_/X _4287_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_100_267 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_619 VGND VPWR sky130_fd_sc_hd__fill_2
X_3238_ _2886_/X _2906_/X _3238_/C _2907_/X _3238_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__4294__B1 _4293_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_340 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_693 VGND VPWR sky130_fd_sc_hd__decap_8
X_3169_ _3021_/X _3035_/X _3055_/X _3014_/Y _3051_/Y _3174_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__2186__A _2183_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_719 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_674 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2914__A _2914_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3729__B _3730_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2633__B _2633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_402 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4551__D _3909_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_571 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3745__A _4474_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_479 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_47 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_378 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3464__B _3437_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_601 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4397__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_144 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4412__RESET_B _2400_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3480__A _3483_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_115 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_502 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_682 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2835__A1 _4318_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_546 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_50 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_83 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3639__B _3637_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2543__B _3806_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4461__D _4523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_222 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3655__A _3660_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_288 VGND VPWR sky130_fd_sc_hd__fill_2
X_2540_ _2532_/X _2539_/X _2540_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_5_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_326 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2771__B1 _4610_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3374__B _3342_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2471_ _2472_/A _2471_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4189__C _4187_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4210_ _2706_/A _2713_/X _4210_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_95_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_446 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_435 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk_i clk_i clkbuf_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_4141_ _4140_/Y _4197_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_95_254 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_619 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2718__B _2718_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4072_ utmi_data_out_o[3] _4072_/B _4072_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3023_ _4356_/Q _3023_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4291__A3 _2533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_493 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_357 VGND VPWR sky130_fd_sc_hd__fill_2
X_3925_ _3925_/A _3924_/X _3925_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4371__D _3664_/Y VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0_clk_i clkbuf_0_clk_i/X clkbuf_2_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_32_571 VGND VPWR sky130_fd_sc_hd__decap_8
X_3856_ _4536_/Q _3844_/X _3856_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_118_632 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3565__A _3555_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2807_ _2691_/A _2666_/X _2805_/X _2806_/Y _2807_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
X_3787_ _2673_/X _3782_/X _3790_/B _2525_/X _3786_/Y _3787_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_118_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_2738_ _2518_/X _2546_/X _2738_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_118_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_315 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2900__C _4421_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3284__B _3283_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4408_ _4408_/D _2865_/C _2405_/X _4410_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2669_ _2669_/A _3717_/A _2691_/B _2669_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_99_582 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_446 VGND VPWR sky130_fd_sc_hd__fill_2
X_4339_ _4339_/D _3306_/A _2487_/X _4430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2909__A _2909_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_78 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_56 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3731__C _3730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_554 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4546__D _3899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2628__B _2624_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4019__B1 utmi_data_out_o[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2644__A _2643_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_538 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_560 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_508 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_593 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3793__A2 _3782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_232 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3475__A _2900_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_247 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_85 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_508 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_clk_i clkbuf_3_3_0_clk_i/A clkbuf_4_5_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_2_431 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_475 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_464 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2819__A _2639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4456__D _2827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_257 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2808__A1 _2636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4412__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_633 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2554__A _2553_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_154 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3369__B _3369_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3710_ _3708_/X _3679_/A _3704_/X _3709_/X _4471_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__4562__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3641_ outport_data_o[6] _3617_/X _3641_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3572_ _3508_/A _3581_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3385__A _2905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_2523_ _4487_/Q _2523_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_646 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4334__RESET_B _2493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_2454_ _2456_/A _2454_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3832__B _3830_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2385_ _2388_/A _2385_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2729__A _3812_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_265 VGND VPWR sky130_fd_sc_hd__decap_4
X_4124_ _4437_/Q _2579_/X _4124_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4366__D _3405_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4055_ _4007_/X _4037_/X _4050_/X _4054_/Y _4055_/X VGND VPWR sky130_fd_sc_hd__a211o_4
Xclkbuf_5_4_0_clk_i clkbuf_5_4_0_clk_i/A _4560_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_3006_ _3005_/Y _3216_/B _3133_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_91_290 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_633 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2464__A _2460_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_696 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3279__B _3278_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_666 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3908_ utmi_data_in_i[7] _3904_/B _3908_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3775__A2 _3673_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3839_ _4529_/Q _3830_/X _3839_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2983__B1 _2982_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2911__B _2911_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_596 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2735__B1 _2520_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2639__A _2638_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_26 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_563 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_585 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_574 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_298 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4435__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3180__D _3179_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_630 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_652 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_663 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2374__A _2339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_482 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_335 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_463 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4585__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_357 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3189__B _3144_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_474 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_390 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2974__B1 _2902_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2821__B _2802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_585 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3636__C _3636_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3933__A _4563_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_627 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_327 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3652__B _3652_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_563 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_70 VGND VPWR sky130_fd_sc_hd__decap_4
X_2170_ _2168_/A _2170_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4027__A1_N _3957_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_599 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_408 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_685 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2284__A _2283_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_633 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_622 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3099__B _3098_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_176 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_165 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4586__RESET_B _2192_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4515__RESET_B _2277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2731__B _2730_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3624_ _4379_/Q _3620_/B _3626_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4004__A _2736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_432 VGND VPWR sky130_fd_sc_hd__fill_2
X_3555_ _3555_/A _3553_/Y _3554_/X _4409_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_3486_ _3516_/A _3486_/B _3486_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3390__B1 _3389_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2506_ _2504_/A _2506_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3562__B _3562_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4458__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_530 VGND VPWR sky130_fd_sc_hd__fill_2
X_2437_ _2434_/A _2437_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2459__A _2456_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_541 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_27_0_clk_i clkbuf_4_13_0_clk_i/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3693__B2 _3692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_2368_ _2367_/X _2368_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_416 VGND VPWR sky130_fd_sc_hd__decap_8
X_2299_ _2301_/A _2299_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4107_ _3964_/A _4039_/B _4033_/A _4106_/Y _4107_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_84_566 VGND VPWR sky130_fd_sc_hd__fill_2
X_4038_ _4030_/X _4039_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2906__B _2905_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2194__A _2188_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_611 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_452 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_149 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2922__A _4330_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_658 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3737__B _3737_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_548 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3175__D _3175_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2369__A _2367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3191__C _3191_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3684__B2 _3669_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_522 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_514 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_633 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_558 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_3_0_clk_i_A clkbuf_5_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_655 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_474 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_72 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2832__A inport_data_i[0] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3928__A _3928_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3647__B _3646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2947__B1 _4428_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_281 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4600__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3663__A _3508_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3340_ _3559_/A _3329_/X _3340_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3372__B1 _3367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_102 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3382__B _3376_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3271_ _3251_/X _3269_/X _3270_/X _4331_/Q _3248_/X _3271_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_112_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_669 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2279__A _2277_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3124__B1 _3014_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4197__C _4199_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_619 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_2222_ _2217_/X _2222_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_23_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_382 VGND VPWR sky130_fd_sc_hd__decap_4
X_2153_ _2155_/A _2153_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_93_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_430 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_282 VGND VPWR sky130_fd_sc_hd__fill_2
X_2986_ _2986_/A _2986_/B _2986_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_30_691 VGND VPWR sky130_fd_sc_hd__fill_2
X_3607_ _3607_/A _3589_/X _3607_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4587_ _4175_/X _4587_/Q _2191_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_115_240 VGND VPWR sky130_fd_sc_hd__decap_4
X_3538_ _3510_/A _3541_/B _3539_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3573__A _2855_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_413 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3292__B _3292_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_295 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_457 VGND VPWR sky130_fd_sc_hd__fill_2
X_3469_ _3498_/A _3528_/D _3528_/A _3528_/B _3486_/B VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_67_39 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2189__A _2188_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3115__B1 _3094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_479 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_680 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2917__A _2917_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_544 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_235 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_38 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_clk_i clkbuf_4_1_0_clk_i/A clkbuf_5_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__4554__D _4554_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_290 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4437__RESET_B _2370_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_87 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3748__A _3749_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_636 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3467__B _3467_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_691 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_64 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_75 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_323 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3483__A _3483_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_566 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4464__D _4526_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2546__B _2546_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_430 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2617__C1 _2616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4082__B2 _4081_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2840_ inport_data_i[4] inport_accept_o _2840_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2967__A1_N _3488_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _4266_/A _4494_/Q _4610_/Q _2770_/Y _2771_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_505 VGND VPWR sky130_fd_sc_hd__fill_2
X_4510_ _4511_/Q _4510_/Q _2283_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4441_ _2723_/X _2707_/A _2365_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_700 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3896__A1 _4545_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4372_ _4303_/X _4372_/Q _2448_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_98_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_3323_ _3317_/A _3322_/X _3323_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4001__B _4000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_3254_ _2917_/A _3266_/B _3254_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_86_628 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_500 VGND VPWR sky130_fd_sc_hd__fill_2
X_2205_ _2206_/A _2205_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_363 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_341 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_566 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_555 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_706 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_717 VGND VPWR sky130_fd_sc_hd__fill_2
X_3185_ _4346_/Q _3186_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_94_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_588 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4374__D _4374_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_547 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_238 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4530__RESET_B _2259_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_377 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_208 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3568__A _3555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2472__A _2472_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2903__C _3464_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2969_ _2926_/A _2965_/A _2968_/Y _2969_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_10_639 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4128__A2 _4127_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_400 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_593 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4549__D _3905_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_433 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_639 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_319 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3750__B _3748_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_650 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2647__A _4527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_330 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4300__A2 _4299_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_160 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4618__RESET_B _2153_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4064__A1 _4562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3682__A1_N _3668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4064__B2 _3933_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3478__A _4420_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2382__A _2396_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3811__A1 _2649_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_591 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_411 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_230 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3697__A1_N _3684_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3925__B _3924_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3878__A1 _4537_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_11_0_clk_i_A clkbuf_4_5_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4459__D _4521_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_552 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4519__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3941__A _4564_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3660__B _3498_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_370 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_469 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_609 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2557__A _2556_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_694 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4359__RESET_B _2463_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_536 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_664 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_193 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_355 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4055__A1 _4007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3388__A _3388_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3941_ _4564_/Q _3941_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_16_282 VGND VPWR sky130_fd_sc_hd__decap_4
X_3872_ _3824_/X _3877_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_90_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2292__A _2288_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2823_ _2796_/A _2818_/X _2822_/X _2823_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_31_285 VGND VPWR sky130_fd_sc_hd__decap_12
X_2754_ _2548_/Y _4282_/B _2753_/X _2754_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_117_324 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4571__SET_B _2211_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2685_ _3717_/A _3713_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3318__B1 _2887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_519 VGND VPWR sky130_fd_sc_hd__decap_12
X_4424_ _4424_/D _3491_/A _2386_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4012__A utmi_data_out_o[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_541 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4369__D _3660_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4355_ _3349_/Y _4355_/Q _2469_/X _4356_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_563 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3851__A _4534_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_628 VGND VPWR sky130_fd_sc_hd__decap_3
X_3306_ _3306_/A _3246_/A _3306_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_58_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3570__B _3582_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4286_ _3808_/A _4498_/Q _4285_/Y _2537_/X _4286_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4294__A1 _3657_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3237_ _4342_/Q _3238_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_39_352 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2467__A _2381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_311 VGND VPWR sky130_fd_sc_hd__decap_4
X_3168_ _3219_/A _3036_/X _3220_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_27_514 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_152 VGND VPWR sky130_fd_sc_hd__fill_1
X_3099_ _3084_/A _3098_/Y _3221_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_14_219 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3298__A _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_79 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_33 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2930__A _2930_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_469 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_44 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_66 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_613 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_403 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3480__B _3478_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_436 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2377__A _2379_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_480 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4452__RESET_B _2352_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2835__A2 _2831_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_558 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_539 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3796__B1 _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3639__C _3639_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2543__C _4502_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_594 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_583 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2840__A inport_data_i[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_296 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3936__A _3186_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3655__B _3653_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2771__B2 _2770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4341__CLK _4430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2470_ _2472_/A _2470_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_79_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_495 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4189__D _4189_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3671__A _3695_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_712 VGND VPWR sky130_fd_sc_hd__decap_12
X_4140_ _4201_/A _4140_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_110_511 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4491__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_469 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2287__A _2283_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4071_ utmi_data_out_o[3] _4072_/B _4071_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_95_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_480 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_171 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_3022_ _4355_/Q _3105_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_64_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_472 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_355 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_580 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3787__B1 _2525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4007__A _4007_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3924_ _2610_/A _3922_/Y _2610_/Y _3923_/Y _3924_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_118_600 VGND VPWR sky130_fd_sc_hd__fill_2
X_3855_ _3883_/A _3855_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2750__A _3814_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2806_ _2638_/Y _2679_/X _2806_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_3786_ _2696_/A _3790_/B _3785_/X _3786_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
Xclkbuf_5_0_0_clk_i clkbuf_5_1_0_clk_i/A _4595_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3565__B _3565_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2737_ _2724_/X _2735_/X _2736_/X _4446_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_118_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_176 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_327 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2900__D _2900_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2668_ _2667_/X _2691_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_4407_ _4407_/D _4407_/Q _2406_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_338 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_319 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3581__A _3581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_561 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_550 VGND VPWR sky130_fd_sc_hd__decap_4
X_2599_ _3994_/A _4437_/Q _2599_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_13 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_200 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_436 VGND VPWR sky130_fd_sc_hd__fill_2
X_4338_ _3305_/Y _3302_/A _2488_/X _4430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_86_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_17 VGND VPWR sky130_fd_sc_hd__fill_1
X_4269_ _4237_/Y _4253_/A _4271_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2197__A _2199_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_288 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2628__C _2628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2925__A _2924_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4019__A1 _4017_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4019__B2 _4018_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4102__A2_N _4108_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_16 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2644__B _4524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3778__B1 _3777_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4562__D _4562_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_32 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_701 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_712 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3793__A3 _3790_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_391 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2660__A _2647_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4364__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_644 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3475__B _3478_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_259 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_299 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3950__B1 _2552_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3491__A _3491_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2819__B _2698_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_704 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_428 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2808__A2 _2803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_461 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_601 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_122 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3218__C1 _3171_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4472__D _4472_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3769__B1 _4472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_133 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3326__A2_N _3325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_572 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3666__A _2826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_391 VGND VPWR sky130_fd_sc_hd__decap_3
X_3640_ _4384_/Q _3640_/B _3642_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_3571_ _3555_/A _3571_/B _3571_/C _3571_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3385__B _2877_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2522_ _4486_/Q _2522_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_53_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_124 VGND VPWR sky130_fd_sc_hd__fill_2
X_2453_ _2425_/A _2456_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_2384_ _2388_/A _2384_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4374__RESET_B _2445_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2729__B _4505_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_564 VGND VPWR sky130_fd_sc_hd__decap_4
X_4123_ _2577_/Y _4122_/X _2608_/Y _4123_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_29_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_406 VGND VPWR sky130_fd_sc_hd__fill_2
X_4054_ _4073_/A _4054_/B _4053_/X _4054_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_110_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_299 VGND VPWR sky130_fd_sc_hd__fill_2
X_3005_ _3005_/A _3005_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_64_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2745__A _4219_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4387__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4382__D _3636_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_678 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_144 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_509 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_19 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3576__A _2855_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3907_ _3889_/A _3897_/X _3906_/X _3907_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_20_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_3838_ _2673_/X _3827_/X _3837_/X _3838_/X VGND VPWR sky130_fd_sc_hd__a21o_4
Xclkbuf_5_23_0_clk_i clkbuf_5_22_0_clk_i/A _4334_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__2983__A1 _3302_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_575 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2480__A _2475_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_708 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_474 VGND VPWR sky130_fd_sc_hd__decap_3
X_3769_ _3680_/Y _3746_/X _4472_/Q _3747_/Y _3769_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2735__A1 _4278_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2735__B2 _2518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3932__B1 _2610_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_56 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4200__A _4198_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_233 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4557__D _4557_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_597 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_620 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2655__A _2680_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_675 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_3_0_clk_i_A clkbuf_4_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_634 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_442 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_431 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_486 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_328 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__A _3516_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_531 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2390__A _2391_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2974__B2 _2973_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_96 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3652__C _3651_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_520 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4475__SET_B _2325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4467__D _4305_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_295 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_534 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_236 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_631 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4100__B1 _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2565__A _4620_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_664 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_420 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_81 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_442 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3396__A _2859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_199 VGND VPWR sky130_fd_sc_hd__decap_4
X_3623_ _3612_/A _3623_/B _3623_/C _3623_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_115_400 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3914__B1 _2571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4004__B _4003_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3554_ _3554_/A _3544_/B _3554_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4555__RESET_B _2229_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_606 VGND VPWR sky130_fd_sc_hd__decap_4
X_3485_ _2900_/D _3478_/B _3485_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3390__A1 _3353_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2505_ _2504_/A _2505_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_639 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3562__C _3561_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_520 VGND VPWR sky130_fd_sc_hd__decap_4
X_2436_ _2434_/A _2436_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4377__D _3655_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_683 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_512 VGND VPWR sky130_fd_sc_hd__decap_3
X_2367_ _2339_/A _2367_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_193 VGND VPWR sky130_fd_sc_hd__fill_1
X_2298_ _2301_/A _2298_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4106_ _4079_/A _4104_/Y _4105_/X _4106_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_84_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2475__A _2496_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4037_ _4079_/A _4037_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_37_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_69 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_667 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_475 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2922__B _2922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3737__C _3736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_394 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3905__B1 _3904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_433 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4402__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_488 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_672 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3191__D _3190_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4552__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_694 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2892__B1 _2867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_214 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2385__A _2388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_589 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_537 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_623 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_283 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2832__B inport_accept_o VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3928__B _2560_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_659 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_9 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2947__B2 _2946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_7_0_clk_i_A clkbuf_4_3_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4105__A _4105_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_219 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3944__A _4321_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_343 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3663__B _3437_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3372__A1 _3337_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3270_ _4331_/Q _3266_/B _3270_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3124__A1 _3227_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_593 VGND VPWR sky130_fd_sc_hd__fill_2
X_2221_ _2217_/X _2221_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_320 VGND VPWR sky130_fd_sc_hd__decap_4
X_2152_ _2252_/A _2155_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_3 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2295__A _2252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_261 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_637 VGND VPWR sky130_fd_sc_hd__decap_4
X_2985_ _2947_/Y _2978_/X _2981_/Y _2984_/Y _2985_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_21_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4425__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3772__A2_N _3771_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3606_ _3415_/Y _3612_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4586_ _4171_/X _4168_/A _2192_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3537_ _4404_/Q _3543_/B _3537_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3573__B _3566_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_615 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4575__CLK _4574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_58 VGND VPWR sky130_fd_sc_hd__decap_3
X_3468_ _3498_/C _3528_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_89_659 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_469 VGND VPWR sky130_fd_sc_hd__fill_1
X_2419_ _2419_/A _2419_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_76_309 VGND VPWR sky130_fd_sc_hd__decap_12
X_3399_ _3399_/A _3399_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_57_501 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3115__B2 _3114_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2917__B _2917_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_383 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_409 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_548 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2933__A _2932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3748__B _3747_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_294 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3467__C _3466_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_456 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4570__D _4570_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2981__A2_N _3298_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4406__RESET_B _2407_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4026__A1_N _4099_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_313 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3483__B _3481_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_285 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4303__B1 _3660_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_158 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_504 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_515 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_206 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2617__B1 _2516_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_261 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3939__A _3939_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4448__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_294 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_283 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_412 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4480__D _3751_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2770_ _4493_/Q _2770_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_8_630 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_681 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_489 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_663 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3674__A _3715_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4440_ _2762_/X _2761_/A _2366_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_7_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_685 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4598__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3896__A2 _3883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_712 VGND VPWR sky130_fd_sc_hd__decap_12
X_4371_ _3664_/Y _3498_/C _2449_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3322_ _2849_/A _3319_/X _3320_/Y _2905_/A _3321_/X _3322_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_3253_ _3253_/A _2956_/X _3253_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_288 VGND VPWR sky130_fd_sc_hd__decap_3
X_2204_ _2206_/A _2204_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3184_ _3181_/X _3183_/Y _4345_/D VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_81_356 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3849__A _4533_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_367 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2753__A _2752_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3568__B _3566_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_434 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2903__D _3653_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4390__D _3605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_445 VGND VPWR sky130_fd_sc_hd__fill_2
X_2968_ _2968_/A _2968_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3584__A _3581_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2899_ _2891_/Y _2892_/Y _2898_/X _2899_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_118_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_412 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2544__C1 _2543_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4569_ _4068_/X _4569_/Q _2213_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_103_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_445 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_327 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_338 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_478 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2928__A _2928_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3750__C _3749_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_117 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_640 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2847__B1 _2846_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4565__D _4565_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_526 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_504 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4049__C1 _4048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_559 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3759__A _3759_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2663__A _2680_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_389 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_710 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4064__A2 _4563_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_209 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3478__B _3478_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3811__A2 _3803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_283 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_242 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_405 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3494__A _3494_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_666 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_644 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3878__A2 _3869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_165 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_58 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_404 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_61 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_106 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2838__A inport_data_i[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_448 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_437 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3660__C _3660_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4475__D _3718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_15_0_clk_i_A clkbuf_4_7_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_673 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_504 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_632 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_345 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_548 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3669__A _3683_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2573__A _2555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4055__A2 _4037_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3940_ _2572_/X _3938_/Y _2611_/X _4043_/A _3940_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3263__B1 _4329_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4399__RESET_B _2415_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4328__RESET_B _2500_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3871_ _4534_/Q _3869_/X _3870_/X _3871_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_83_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2822_ _2691_/A _2820_/X _2624_/A _2821_/Y _2822_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_31_264 VGND VPWR sky130_fd_sc_hd__decap_4
X_2753_ _2752_/X _2753_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_336 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3318__A1 _4376_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2684_ _2669_/A _2684_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4423_ _4423_/D _3488_/A _2387_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4354_ _3339_/Y _4354_/Q _2470_/X _4356_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_575 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3851__B _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_607 VGND VPWR sky130_fd_sc_hd__decap_3
X_3305_ _3317_/A _3304_/Y _3305_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2748__A _4499_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4285_ _4502_/Q _3816_/A _4506_/Q _4285_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_104_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_459 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4385__D _3645_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3236_ _3366_/A _3235_/X _3236_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4294__A2 _4292_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4613__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3757__A1_N _3683_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_59 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_470 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3127__A1_N _3050_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3167_ _3205_/C _3088_/Y _3166_/X _3167_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_81_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_345 VGND VPWR sky130_fd_sc_hd__fill_2
X_3098_ _3097_/X _3098_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_120_14 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3579__A _4400_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_507 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2483__A _2485_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3298__B _3298_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_570 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2930__B _2948_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_303 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_78 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_89 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2658__A _4525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3480__C _3480_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_597 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_407 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_18_0_clk_i clkbuf_4_9_0_clk_i/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_651 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_429 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_632 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2393__A _2391_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3489__A _3547_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_687 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_518 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4492__RESET_B _2305_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_581 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4421__RESET_B _2390_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3796__A1 _2684_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3796__B2 _3792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_231 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2543__D _4503_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3936__B _4278_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2840__B inport_accept_o VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_279 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3655__C _3654_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_317 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_463 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3952__A _4322_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2568__A _2580_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_691 VGND VPWR sky130_fd_sc_hd__decap_12
X_4070_ _4012_/Y _4069_/X _4012_/Y _4069_/X _4072_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_92 VGND VPWR sky130_fd_sc_hd__fill_1
X_3021_ _3071_/A _3021_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_76_492 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4509__RESET_B _2284_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3399__A _3399_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_507 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3787__A1 _2673_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3787__B2 _3786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3923_ _4570_/Q _3923_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_551 VGND VPWR sky130_fd_sc_hd__fill_2
X_3854_ _4527_/Q _3841_/X _3853_/X _3854_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_2805_ _2785_/C _2804_/X _2635_/A _2805_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3785_ _3785_/A _3785_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2750__B _3816_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3565__C _3564_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2736_ _2696_/A _2736_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_105_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_2667_ _2785_/C _2666_/X _2667_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4406_ _3545_/Y _3543_/A _2407_/X _4410_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3681__A1_N _3680_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3581__B _3579_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2598_ _3980_/B _3993_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_523 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_415 VGND VPWR sky130_fd_sc_hd__fill_2
X_4337_ _3300_/Y _3297_/A _2490_/X _4334_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2478__A _2475_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_245 VGND VPWR sky130_fd_sc_hd__decap_4
X_4268_ _4265_/A _4266_/X _4267_/Y _4268_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_86_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_470 VGND VPWR sky130_fd_sc_hd__fill_2
X_3219_ _3219_/A _3026_/X _3219_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4199_ _4198_/Y _4199_/B _4199_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_3_3_0_clk_i_A clkbuf_3_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4019__A2 utmi_data_out_o[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_304 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3102__A _3007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3778__A1 _3698_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_11 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4509__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2941__A _2941_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_370 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_724 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_77 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_144 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3950__B2 _3949_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3950__A1 _2578_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3491__B _3479_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_372 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2388__A _2388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_256 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_716 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_237 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4602__RESET_B _2173_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_624 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4108__A _4009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3218__B1 _3217_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3012__A _3007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3769__B2 _3747_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3769__A1 _3680_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_178 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2851__A _2850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3947__A _3947_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_83 VGND VPWR sky130_fd_sc_hd__fill_2
X_3570_ _3513_/A _3582_/B _3571_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3385__C _3332_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_604 VGND VPWR sky130_fd_sc_hd__fill_2
X_2521_ _4228_/B _2724_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_5_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_158 VGND VPWR sky130_fd_sc_hd__decap_12
X_2452_ _2449_/A _2452_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_46_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_2383_ _2388_/A _2383_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_713 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2298__A _2301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_180 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_320 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_223 VGND VPWR sky130_fd_sc_hd__decap_3
X_4122_ _2605_/X _2579_/X _4122_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_418 VGND VPWR sky130_fd_sc_hd__fill_2
X_4053_ utmi_data_out_o[0] _4053_/B _4053_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_83_237 VGND VPWR sky130_fd_sc_hd__decap_3
X_3004_ _2999_/X _3003_/X _2996_/A _3004_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_52_602 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_676 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4343__RESET_B _2483_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2745__B _2548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_484 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4018__A utmi_data_out_o[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_3906_ utmi_data_in_i[6] _3904_/B _3906_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_51_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_156 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2761__A _2761_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3576__B _3566_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_381 VGND VPWR sky130_fd_sc_hd__fill_1
X_3837_ _3837_/A _3830_/X _3837_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2983__A2 _2979_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3768_ _3724_/A _3674_/B _2687_/X _3767_/Y _3768_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_106_615 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2735__A2 _2734_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2719_ _2719_/A _4278_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_4_10_0_clk_i_A clkbuf_3_5_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_208 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3932__A1 _2571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3932__B2 _4041_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3699_ _3683_/Y _3698_/A _3683_/A _3698_/Y _3699_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_105_103 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3592__A outport_data_o[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_629 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_681 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4200__B _4199_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2936__A _3297_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_610 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2655__B _2654_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4331__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_281 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4573__D _4092_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_454 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_134 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7_0_clk_i_A clkbuf_4_7_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3767__A _3708_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2671__A _2671_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4481__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__B _3486_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_420 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_241 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3007__A _4361_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_83 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2846__A inport_data_i[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4100__B2 _4022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2565__B _3994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_654 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4483__D _3768_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_454 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_93 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3677__A _3677_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_370 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2581__A _2581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3396__B _3398_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3622_ outport_data_o[0] _3625_/B _3623_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_412 VGND VPWR sky130_fd_sc_hd__decap_8
X_3553_ _2865_/B _3541_/B _3553_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3914__B2 _4569_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_467 VGND VPWR sky130_fd_sc_hd__fill_2
X_3484_ _3660_/A _3504_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3390__A2 _3394_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2504_ _2504_/A _2504_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_478 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_117 VGND VPWR sky130_fd_sc_hd__decap_4
X_2435_ _2434_/A _2435_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4595__RESET_B _2182_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_351 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4524__RESET_B _2266_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2366_ _2362_/A _2366_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4105_ _4105_/A _4103_/X _4105_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_84_546 VGND VPWR sky130_fd_sc_hd__fill_2
X_2297_ _2301_/A _2297_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4354__CLK _4356_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_4036_ _4030_/X _4079_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4393__D _4393_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_602 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3850__B1 _3849_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3587__A _3586_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_129 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2491__A _2495_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_329 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3905__A1 _4549_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4481__SET_B _2318_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_528 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_456 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4211__A _3987_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4568__D _4063_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_437 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4241__A1_N _4242_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2666__A _4450_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2892__B2 _2874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2892__A1 _2877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_101 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_97 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_646 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3497__A _3428_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_616 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4105__B _4103_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_322 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_250 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3944__B _3944_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_399 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3372__A2 _3371_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4121__A _2566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4478__D _3738_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4377__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3960__A _4323_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3124__A2 _3080_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2220_ _2217_/X _2220_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_78_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_535 VGND VPWR sky130_fd_sc_hd__fill_2
X_2151_ _2381_/A _2252_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2576__A _2572_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_527 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_605 VGND VPWR sky130_fd_sc_hd__fill_2
X_2984_ _3451_/A _3303_/B _3451_/A _3303_/B _2984_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_15_690 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3899__B1 _3898_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3605_ _3585_/X _3603_/X _3604_/X _3605_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4585_ _4585_/D _4585_/Q _2193_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3536_ _3545_/A _3534_/Y _3536_/C _4403_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4031__A _4010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_627 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4388__D _3599_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3870__A _4542_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3467_ _3483_/A _3467_/B _3466_/X _3467_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_97_660 VGND VPWR sky130_fd_sc_hd__fill_2
X_2418_ _2419_/A _2418_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3398_ _2859_/A _3398_/B _3398_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_96_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_310 VGND VPWR sky130_fd_sc_hd__fill_2
X_2349_ _2352_/A _2349_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2486__A _2485_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_387 VGND VPWR sky130_fd_sc_hd__decap_8
X_4019_ _4017_/Y utmi_data_out_o[4] utmi_data_out_o[0] _4018_/Y _4019_/X VGND VPWR
+ sky130_fd_sc_hd__o22a_4
XANTENNA__4076__B1 _4011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_454 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_593 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_284 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_649 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_487 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4206__A _4205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3110__A _3011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_592 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4008__A2_N _4007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4000__B1 _3962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3483__C _3483_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4446__RESET_B _2359_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2562__B1 _2908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4303__A1 _4372_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3780__A _3707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2396__A _2396_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_470 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_535 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_524 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_527 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2617__A1 _2595_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_443 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_465 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_593 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4116__A _4116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_424 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3020__A _4354_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3955__A _3955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_660 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_653 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3674__B _3674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_174 VGND VPWR sky130_fd_sc_hd__fill_2
X_4370_ _3662_/X _3528_/C _2450_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_3321_ _3234_/Y _2992_/Y _3319_/A _3244_/B _3321_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_112_223 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3690__A _3690_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_435 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_424 VGND VPWR sky130_fd_sc_hd__decap_4
X_3252_ _3265_/A _3253_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_79_660 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_310 VGND VPWR sky130_fd_sc_hd__decap_12
X_2203_ _2206_/A _2203_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3183_ _3928_/A _2999_/X _3240_/A _3183_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_93_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_579 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4058__B1 _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3849__B _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_560 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3568__C _3567_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3865__A _4540_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2967_ _3488_/A _2966_/X _3488_/A _2966_/X _2967_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_10_619 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_479 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4542__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2898_ _2896_/X _2897_/Y _2898_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_118_14 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3584__B _3582_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2792__B1 _2636_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2544__B1 _2540_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4568_ _4063_/X _4568_/Q _2214_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_1_306 VGND VPWR sky130_fd_sc_hd__decap_6
X_3519_ _3547_/A _3516_/B _3520_/C VGND VPWR sky130_fd_sc_hd__and2_4
X_4499_ _3809_/Y _4499_/Q _2297_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_103_245 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2928__B _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4297__B1 _2684_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_129 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2847__A1 _4324_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3105__A _3015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4049__B1 _4033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_538 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_66 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3759__B _3770_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2663__B _2662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_722 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4581__D _4151_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_428 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4221__B1 _2704_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_14_0_clk_i clkbuf_4_7_0_clk_i/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3494__B _3479_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_634 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_133 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_521 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3732__C1 _3731_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2838__B inport_accept_o VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_416 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_350 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3015__A _4356_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4415__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_655 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_644 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_72 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2854__A _2854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3263__A1 _3251_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3669__B _4474_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_19_0_clk_i_A clkbuf_4_9_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_508 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_700 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3263__B2 _3248_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_176 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4491__D _4491_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3870_ _4542_/Q _3859_/B _3870_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3156__A2_N _3070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4565__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_232 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3685__A _4522_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2821_ _2821_/A _2802_/X _2821_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_76_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_2752_ _4278_/D _2761_/C _2752_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2774__B1 _4236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4368__RESET_B _2452_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_359 VGND VPWR sky130_fd_sc_hd__decap_3
X_4422_ _4422_/D _2900_/D _2388_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2683_ _2671_/A _2631_/X _2682_/X _2681_/Y _2683_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3318__A2 _2906_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4087__A1_N _3957_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4353_ _2890_/Y _4353_/Q _2471_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_101_705 VGND VPWR sky130_fd_sc_hd__fill_2
X_3304_ _3280_/X _3302_/X _3303_/X _3302_/A _3248_/A _3304_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_4284_ _2533_/X _4283_/B _2548_/A _4284_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4010__A1_N _4008_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_298 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_3235_ _3319_/A _3234_/Y _3244_/B _3235_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__2748__B _4498_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_clk_i_A clkbuf_2_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_663 VGND VPWR sky130_fd_sc_hd__fill_2
X_3166_ _3070_/X _3363_/A _3061_/X _3110_/C _3166_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_81_110 VGND VPWR sky130_fd_sc_hd__fill_2
X_3097_ _3031_/X _3347_/B _3359_/A _3359_/B _3097_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3579__B _3582_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_593 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_582 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_390 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_541 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_563 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4203__B1 _4143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_3999_ _4602_/Q _3999_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3595__A outport_data_o[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_39 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_392 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3714__C1 _3713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2939__A _2938_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_254 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4576__D _4576_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4438__CLK _4574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_630 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_460 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_674 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2674__A _4524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_622 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3489__B _3486_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_655 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_154 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4588__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_305 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_700 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3796__A2 _3785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4461__RESET_B _2342_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2756__B1 _2602_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2849__A _2849_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3952__B _2585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4486__D _4486_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_427 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2568__B _2568_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_685 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_140 VGND VPWR sky130_fd_sc_hd__decap_3
X_3020_ _4354_/Q _3071_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_5_30_0_clk_i_A clkbuf_5_30_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2584__A _3944_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_699 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4549__RESET_B _2236_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3787__A2 _3782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_198 VGND VPWR sky130_fd_sc_hd__fill_2
X_3922_ _2604_/X _3919_/Y _3920_/X _2581_/A _3921_/Y _3922_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_3853_ _4535_/Q _3844_/X _3853_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_703 VGND VPWR sky130_fd_sc_hd__decap_4
X_2804_ _2804_/A _3704_/A _2804_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4304__A _2639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_101 VGND VPWR sky130_fd_sc_hd__decap_4
X_3784_ _3784_/A _3790_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2750__C _2750_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_646 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_123 VGND VPWR sky130_fd_sc_hd__fill_2
X_2735_ _4278_/D _2734_/X _2520_/Y _2518_/X _2735_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_8_280 VGND VPWR sky130_fd_sc_hd__decap_12
X_2666_ _4450_/Q _2666_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4405_ _3542_/Y _4405_/Q _2408_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_530 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2759__A _4468_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3581__C _3581_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4336_ _3296_/Y _3293_/A _2491_/X _4334_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2597_ _3994_/B _3980_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4396__D _3568_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_405 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_48 VGND VPWR sky130_fd_sc_hd__fill_2
X_4267_ _4267_/A _4264_/B _4267_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_55_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_600 VGND VPWR sky130_fd_sc_hd__fill_2
X_3218_ _3019_/Y _3085_/B _3217_/Y _3171_/B _3218_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_4198_ _4592_/Q _4198_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2494__A _2495_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_493 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_644 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_3149_ _3073_/Y _3114_/X _3153_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_655 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_508 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_636 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_316 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3102__B _3038_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_379 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3778__A2 _3776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_i_A clkbuf_3_7_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_390 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_23 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_382 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_585 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3950__A2 _3948_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2669__A _2669_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3163__B1 _3240_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_202 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_489 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3173__A1_N _3041_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_224 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_357 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4108__B _4108_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3218__A1 _3019_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3769__A2 _3746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_658 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_338 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3012__B _3008_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2977__B1 _4427_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4124__A _4437_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3385__D _2872_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4603__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2520_ _4446_/Q _2520_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2451_ _2449_/A _2451_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2579__A _2578_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3154__B1 _3085_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_500 VGND VPWR sky130_fd_sc_hd__fill_2
X_2382_ _2396_/A _2388_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_533 VGND VPWR sky130_fd_sc_hd__decap_4
X_4121_ _2566_/X _4120_/Y _4127_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4052_ utmi_data_out_o[0] _4053_/B _4054_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_110_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_216 VGND VPWR sky130_fd_sc_hd__decap_12
X_3003_ _3003_/A _3248_/A _3003_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_37_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_430 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2745__C _4469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3203__A _2996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_496 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_614 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_699 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_688 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_293 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2950__A1_N _3494_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_658 VGND VPWR sky130_fd_sc_hd__decap_8
X_3905_ _4549_/Q _3897_/X _3904_/X _3905_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4383__RESET_B _2435_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2761__B _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_393 VGND VPWR sky130_fd_sc_hd__decap_4
X_3836_ utmi_rxvalid_i _4519_/Q utmi_rxactive_i _4519_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4034__A _4561_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_544 VGND VPWR sky130_fd_sc_hd__decap_12
X_3767_ _3708_/A _3765_/X _3766_/Y _3767_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_118_454 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3873__A _4543_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3393__B1 _3392_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2718_ _2716_/Y _2718_/B _2719_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3932__A2 _3930_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3698_ _3698_/A _3698_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_498 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_115 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3592__B _3592_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_148 VGND VPWR sky130_fd_sc_hd__fill_2
X_2649_ _4522_/Q _2649_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2489__A _2496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_619 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3696__A1 _3671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14_0_clk_i_A clkbuf_3_7_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_213 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_544 VGND VPWR sky130_fd_sc_hd__fill_1
X_4319_ _2837_/X _4319_/Q _2510_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_75_706 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2936__B _2935_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3113__A _3048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_688 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_349 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2959__B1 _2958_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3767__B _3765_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_308 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2671__B _2669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_360 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_32 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_526 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3783__A _2624_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_476 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2399__A _2399_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3136__B1 _3066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_253 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_555 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_685 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2846__B _2846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_569 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_709 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3023__A _4356_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4119__A _3993_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_614 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_699 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2862__A _2862_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_61 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_647 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2764__A2_N _4496_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_466 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3677__B _3676_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_680 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_382 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_218 VGND VPWR sky130_fd_sc_hd__fill_2
X_3621_ _3617_/X _3625_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_3552_ _3555_/A _3550_/Y _3552_/C _4408_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_2503_ _2496_/A _2504_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_581 VGND VPWR sky130_fd_sc_hd__fill_2
X_3483_ _3483_/A _3481_/Y _3483_/C _4421_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_6_592 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3127__B1 _3045_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2434_ _2434_/A _2434_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_500 VGND VPWR sky130_fd_sc_hd__fill_2
X_2365_ _2362_/A _2365_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_706 VGND VPWR sky130_fd_sc_hd__decap_12
X_4104_ _4105_/A _4103_/X _4104_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_110_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_2296_ _2324_/A _2301_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_37_452 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4029__A _3994_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4035_ _4561_/Q _4034_/B _4033_/X _4034_/Y _4561_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_112_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_474 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_102 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3850__A1 _4525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_591 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_636 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_119 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_319 VGND VPWR sky130_fd_sc_hd__fill_2
X_3819_ _2650_/Y _3804_/B _3818_/X _4504_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_4_507 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3905__A2 _3897_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_7 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_68 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_446 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_28 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4211__B _2704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3118__B1 _3219_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3108__A _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_449 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_396 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2892__A2 _2872_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4584__D _4163_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_506 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_260 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4238__A2_N _4260_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_591 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2682__A _2669_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_135 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_477 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_455 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_64 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_691 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_138 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_352 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3357__B1 _3356_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4121__B _4120_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3109__B1 _3381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_540 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3018__A _3017_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3960__B _3960_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_72 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2857__A _2857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_482 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_514 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2576__B _2575_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2150_ rst_i _2381_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4494__D _3798_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_377 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_506 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_274 VGND VPWR sky130_fd_sc_hd__fill_2
X_2983_ _3302_/A _2979_/A _2982_/Y _3303_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_14_190 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3348__B1 _3366_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3899__A1 _4546_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3604_ outport_data_o[4] _3592_/B _3604_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4584_ _4163_/X _4160_/A _2194_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3535_ _3506_/A _3541_/B _3536_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4031__B _4031_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_639 VGND VPWR sky130_fd_sc_hd__decap_12
X_3466_ _3554_/A _3462_/B _3466_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4321__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_287 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3870__B _3859_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2417_ _2396_/A _2419_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_127 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_341 VGND VPWR sky130_fd_sc_hd__decap_12
X_3397_ _3397_/A _3394_/Y _3396_/Y _4364_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_97_672 VGND VPWR sky130_fd_sc_hd__decap_6
X_2348_ _2352_/A _2348_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_536 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4471__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_493 VGND VPWR sky130_fd_sc_hd__fill_1
X_2279_ _2277_/A _2279_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_558 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_219 VGND VPWR sky130_fd_sc_hd__fill_2
X_4018_ utmi_data_out_o[4] _4018_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4076__B2 _4075_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3598__A outport_data_o[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_13 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_477 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3110__B _3369_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_56 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3339__B1 _3338_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_711 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4222__A _4116_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4000__A1 _3999_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4000__B2 _3981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4579__D _4142_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2562__A1 inport_valid_i VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2562__B2 _4278_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_359 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3780__B _3780_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_521 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_108 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2677__A _2676_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4303__A2 _3420_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4486__RESET_B _2312_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_53 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4415__RESET_B _2397_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_10_0_clk_i clkbuf_4_5_0_clk_i/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_87_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_355 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_539 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2617__A2 _4033_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3301__A _3240_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_85 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4100__A2_N _4022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_488 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4116__B _3984_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_458 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_469 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_672 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_7 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3674__C _3674_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_142 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4132__A _3993_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4344__CLK _4325_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4489__D _4489_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_414 VGND VPWR sky130_fd_sc_hd__fill_1
X_3320_ _3653_/A _3320_/B _3320_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3971__A _3229_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_82 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4494__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_469 VGND VPWR sky130_fd_sc_hd__fill_2
X_3251_ _3251_/A _3251_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_94_620 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_171 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_514 VGND VPWR sky130_fd_sc_hd__fill_2
X_2202_ _2166_/X _2206_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_21_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_3182_ _3182_/A _3928_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_94_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_322 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_675 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4058__B2 _3925_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_293 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3211__A _3392_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_252 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4307__A _2706_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_2966_ _4331_/Q _2951_/A _2965_/Y _2966_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3865__B _3859_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2897_ _4379_/Q _2880_/A _3331_/D _2876_/A _2872_/B _2897_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
XFILLER_30_491 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3584__C _3583_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2792__A1 _2804_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4399__D _4399_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_552 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3881__A _4547_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3741__B1 _3708_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_19 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2544__A1 _2534_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4567_ _4055_/X _4007_/A _2215_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_116_585 VGND VPWR sky130_fd_sc_hd__decap_8
X_3518_ _2864_/D _3512_/B _3518_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_89_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_4498_ _3807_/Y _4498_/Q _2298_/X _4450_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2497__A _2497_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3449_ _3513_/A _3462_/B _3449_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4297__A1 _2528_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2847__A2 _2829_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3105__B _4357_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4049__A1 _4566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_358 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_583 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_11 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3121__A _3120_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_403 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4367__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_458 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_296 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4208__A1_N _4207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_255 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4221__A1 _4595_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4221__B2 _2755_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_480 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_563 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3732__B1 _3719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3791__A _3785_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3167__B1_N _3166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2200__A _2199_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_395 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_539 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3669__C _3669_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3799__B1 _4525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4127__A _2612_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3263__A2 _3261_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_188 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_263 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3031__A _4354_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_200 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3966__A _4007_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2820_ _2636_/A _2819_/Y _2785_/X _2820_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__2870__A _3331_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2751_ _2711_/X _2750_/X _2761_/C VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_491 VGND VPWR sky130_fd_sc_hd__fill_2
X_2682_ _2669_/A _3717_/A _2666_/X _2682_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__2774__B2 _2773_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4421_ _4421_/D _4421_/Q _2390_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_69_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4069__A2_N _4022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_222 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4337__RESET_B _2490_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4352_ _2996_/Y _4352_/Q _2472_/X _4325_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3303_ _3253_/A _3303_/B _3303_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4283_ _2533_/X _4283_/B _4283_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_98_288 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_266 VGND VPWR sky130_fd_sc_hd__fill_2
X_3234_ _2913_/B _3234_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3206__A _3350_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_344 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_311 VGND VPWR sky130_fd_sc_hd__fill_2
X_3165_ _3108_/X _3153_/A _3165_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_27_506 VGND VPWR sky130_fd_sc_hd__fill_2
X_3096_ _3227_/D _3094_/X _3095_/X _3112_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_27_528 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_678 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4037__A _4079_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2780__A _2696_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_553 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4203__A1 _2516_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3998_ _3996_/X _3997_/X _2602_/X _4558_/D VGND VPWR sky130_fd_sc_hd__o21a_4
X_2949_ _2928_/A _2968_/A _2948_/Y _2949_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3595__B _3592_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_299 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_327 VGND VPWR sky130_fd_sc_hd__decap_8
X_4619_ _4619_/D _2526_/C _2155_/A _4619_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3714__B1 _3704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_533 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3116__A _3021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_99 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_133 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_10 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_347 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4592__D _4592_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_54 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_572 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3796__A3 _4492_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2690__A _3707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_42 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2756__A1 _2743_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_51 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4430__RESET_B _2378_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_203 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3026__A _3021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_631 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_620 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2865__A _3543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4130__B1 _4231_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4532__CLK _4539_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_420 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_472 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_163 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_358 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_317 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_550 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3787__A3 _3790_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_391 VGND VPWR sky130_fd_sc_hd__fill_2
X_3921_ _4554_/Q _3921_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_542 VGND VPWR sky130_fd_sc_hd__fill_2
X_3852_ _2659_/X _3841_/X _3851_/X _3852_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__2995__A1 _2916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2803_ _2803_/A _2802_/X _2803_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_586 VGND VPWR sky130_fd_sc_hd__fill_2
X_3783_ _2624_/A _2666_/X _3784_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4304__B _2800_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2750__D _2749_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4589__RESET_B _2189_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_113 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4518__RESET_B _2273_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2734_ _2727_/X _2730_/X _2731_/X _4215_/B _2734_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_117_168 VGND VPWR sky130_fd_sc_hd__fill_2
X_2665_ _2671_/A _2631_/X _2664_/X _2671_/D _2665_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_8_292 VGND VPWR sky130_fd_sc_hd__decap_3
X_4404_ _4404_/D _4404_/Q _2409_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_319 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2759__B _2548_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2596_ _2596_/A _3994_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_341 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_542 VGND VPWR sky130_fd_sc_hd__decap_6
X_4335_ _3292_/Y _3289_/A _2492_/X _4334_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_586 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_558 VGND VPWR sky130_fd_sc_hd__fill_2
X_4266_ _4266_/A _4263_/B _4266_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_74_409 VGND VPWR sky130_fd_sc_hd__decap_12
X_3217_ _3146_/X _3217_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4197_ _4197_/A _4197_/B _4199_/B _4197_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_3148_ _3148_/A _3143_/Y _3108_/X _3228_/A _3148_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_27_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_133 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_486 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_615 VGND VPWR sky130_fd_sc_hd__decap_12
X_3079_ _3350_/C _4357_/Q _4354_/Q _4355_/Q _3079_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_70_659 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3102__C _4358_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_520 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_564 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_575 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_636 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_23 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4405__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_680 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_179 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4230__A _4247_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_341 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2669__B _3717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_435 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4587__D _4175_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3163__A1 _3920_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_214 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4555__CLK _4619_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2685__A _3717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_601 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4112__B1 _4030_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_306 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3218__A2 _3085_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3012__C _3010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_520 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2977__B2 _2976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_553 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_586 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4124__B _2579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3926__B1 _3925_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4611__RESET_B _2162_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2450_ _2449_/A _2450_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4140__A _4201_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4497__D _2780_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3154__A1 _3059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_512 VGND VPWR sky130_fd_sc_hd__decap_3
X_2381_ _2381_/A _2396_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_704 VGND VPWR sky130_fd_sc_hd__fill_2
X_4120_ _2579_/X _2572_/X _2575_/X _4120_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_96_589 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_601 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4103__B1 _4100_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4051_ _4561_/Q _3964_/A _3915_/Y _3964_/Y _4053_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2595__A _2595_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_377 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_228 VGND VPWR sky130_fd_sc_hd__fill_2
X_3002_ _3277_/A _3248_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_64_420 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3203__B _3195_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_136 VGND VPWR sky130_fd_sc_hd__fill_2
X_3904_ utmi_data_in_i[5] _3904_/B _3904_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4315__A enable_i VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3090__B1 _3085_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2761__C _2761_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3835_ _4518_/Q _3827_/X _3834_/X _4518_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4428__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4034__B _4034_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_556 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_433 VGND VPWR sky130_fd_sc_hd__fill_2
X_3766_ _3762_/Y _3764_/X _3766_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2947__A2_N _2946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4352__RESET_B _2472_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3873__B _3877_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3393__A1 _3342_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2717_ _2761_/A _2718_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3697_ _3684_/X _3696_/X _3684_/X _3696_/X _3698_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_628 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4578__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_37 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4050__A _4050_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2648_ _4523_/Q _4527_/Q _2648_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_10_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_108 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3696__A2 _3695_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_650 VGND VPWR sky130_fd_sc_hd__fill_1
X_2579_ _2578_/X _2579_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_225 VGND VPWR sky130_fd_sc_hd__fill_2
X_4318_ _2835_/X _4318_/Q _2511_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4249_ _4249_/A _4249_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_101_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_634 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2656__B1 _2655_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3113__B _3098_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_667 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_12 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_177 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_659 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_56 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_188 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2959__A1 _4328_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3767__C _3766_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_478 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_158 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2671__C _2670_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_681 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_512 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_394 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_433 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3783__B _2666_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_609 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_108 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3136__B2 _3045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_287 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_567 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_74 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_431 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4119__B _4118_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_475 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2862__B _4405_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_272 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_478 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4135__A _2669_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_692 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3974__A _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3620_ _4378_/Q _3620_/B _3623_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_3551_ _3522_/A _3544_/B _3552_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_2502_ _2497_/A _2502_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_458 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_436 VGND VPWR sky130_fd_sc_hd__decap_3
X_3482_ _3513_/A _3479_/B _3483_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_51_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_108 VGND VPWR sky130_fd_sc_hd__fill_2
X_2433_ _2434_/A _2433_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3127__B2 _3223_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_545 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2886__B1 _2896_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2364_ _2362_/A _2364_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_504 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_718 VGND VPWR sky130_fd_sc_hd__decap_6
X_4103_ _4100_/X _4102_/X _4100_/X _4102_/X _4103_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_375 VGND VPWR sky130_fd_sc_hd__decap_12
X_2295_ _2252_/A _2324_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3214__A _3367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4029__B _2581_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4034_ _4561_/Q _4034_/B _4034_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_37_464 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_615 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3850__A2 _3841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_114 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_158 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4533__RESET_B _2256_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_692 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_681 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4045__A _4030_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3884__A _3884_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3818_ _3818_/A _3804_/Y _3818_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_230 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_36 VGND VPWR sky130_fd_sc_hd__fill_2
X_3749_ _3749_/A _3747_/Y _3749_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_118_285 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_7 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3118__A1 _3098_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_714 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3108__B _3065_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_491 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_642 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_331 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_675 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_537 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_526 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2892__A3 _2872_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_55 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_272 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_412 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_659 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_72 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2682__B _3717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_242 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_147 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_83 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_489 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_128 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_98 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_375 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3357__A1 _2851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_38 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3109__A1 _3046_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2203__A _2206_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_106 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3109__B2 _3008_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_574 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2857__B _3559_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_718 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_707 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_472 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3034__A _3120_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_367 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2873__A _2872_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3969__A _4568_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_220 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_286 VGND VPWR sky130_fd_sc_hd__fill_2
X_2982_ _2940_/B _2982_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_22_618 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_297 VGND VPWR sky130_fd_sc_hd__decap_4
X_3603_ _2858_/B _3589_/X _3603_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3348__A1 _3346_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_684 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_695 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3899__A2 _3897_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4583_ _4583_/D _4156_/A _2196_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3209__A _3209_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_222 VGND VPWR sky130_fd_sc_hd__fill_2
X_3534_ _4403_/Q _3543_/B _3534_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_266 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_618 VGND VPWR sky130_fd_sc_hd__fill_2
X_3465_ outport_data_o[7] _3554_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2416_ _2411_/A _2416_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_103_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_353 VGND VPWR sky130_fd_sc_hd__decap_12
X_3396_ _2859_/B _3398_/B _3396_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4616__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_472 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_461 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_301 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_375 VGND VPWR sky130_fd_sc_hd__fill_1
X_2347_ _2352_/A _2347_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_526 VGND VPWR sky130_fd_sc_hd__fill_2
X_2278_ _2277_/A _2278_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_397 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3879__A _4546_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_356 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2783__A _2782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_250 VGND VPWR sky130_fd_sc_hd__fill_2
X_4017_ utmi_data_out_o[0] _4017_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3598__B _3592_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_570 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_25 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_401 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_629 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_448 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3110__C _3110_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_662 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3339__A1 _2851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_723 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3119__A _3119_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_194 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4222__B _4207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4000__A2 _3994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_327 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2958__A _2920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2562__A2 _2557_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_214 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4126__B1_N _2569_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_533 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4595__D _4212_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_450 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3694__A1_N _3687_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_337 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4455__RESET_B _2349_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_42 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_404 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4116__C _4116_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_150 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_509 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3674__D _3674_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_154 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4132__B _4131_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_699 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3029__A _3028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_61 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2868__A _4378_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3971__B _4278_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_3250_ _3268_/A _3249_/Y _3250_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_79_640 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_504 VGND VPWR sky130_fd_sc_hd__decap_4
X_2201_ _2199_/A _2201_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3181_ _3181_/A _3181_/B _3216_/B _3180_/X _3181_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_93_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_209 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_2965_ _2965_/A _2965_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2896_ _2896_/A _4375_/Q _2895_/X _2896_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__2792__A2 _2691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_531 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_4566_ _4049_/X _4566_/Q _2216_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3517_ _3514_/A _3517_/B _3517_/C _4414_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3881__B _3877_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3741__A1 _3680_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2544__A2 _2537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_437 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2778__A _2777_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4497_ _2780_/X _4497_/Q _2299_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_103_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_448 VGND VPWR sky130_fd_sc_hd__decap_12
X_3448_ outport_data_o[3] _3513_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4297__A2 _3960_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3379_ _3317_/A _3379_/B _4360_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_97_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_312 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3105__C _4354_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_518 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4049__A2 _4037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3402__A _2858_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_415 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4221__A2 _2743_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_102 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_542 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3732__A1 _3726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_658 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2688__A _2673_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_64 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_385 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_665 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_52 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3669__D _3668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3799__A1 _2601_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3799__B2 _3792_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4127__B _4127_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_592 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3263__A3 _3262_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_286 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_212 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_2750_ _3814_/A _3816_/A _2750_/C _2749_/X _2750_/X VGND VPWR sky130_fd_sc_hd__or4_4
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4143__A _4140_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4461__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2681_ _3780_/B _2629_/X _2680_/X _2681_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_117_328 VGND VPWR sky130_fd_sc_hd__fill_1
X_4420_ _4420_/D _4420_/Q _2391_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_523 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_4351_ _3004_/Y _4231_/C _2473_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2598__A _3980_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_234 VGND VPWR sky130_fd_sc_hd__fill_2
X_3302_ _3302_/A _3246_/A _3302_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4282_ _4282_/A _4282_/B _2713_/X _2546_/B _4283_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_113_567 VGND VPWR sky130_fd_sc_hd__fill_1
X_3233_ _3231_/Y _3232_/X _3233_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3206__B _3359_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4377__RESET_B _2442_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_356 VGND VPWR sky130_fd_sc_hd__fill_2
X_3164_ _3160_/X _3163_/Y _4344_/D VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_82_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_378 VGND VPWR sky130_fd_sc_hd__decap_12
X_3095_ _3048_/Y _3095_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3222__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_562 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_532 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_223 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2780__B _2779_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_407 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4203__A2 _4202_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3997_ _3994_/A _3994_/B _4558_/Q _3997_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_2948_ _2948_/A _2948_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4053__A utmi_data_out_o[0] VGND VPWR sky130_fd_sc_hd__diode_2
X_2879_ _2876_/A _4379_/Q _2879_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4618_ _4618_/D _2528_/C _2153_/X _4619_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3714__A1 _3708_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4549_ _3905_/X _4549_/Q _2236_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_8 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_617 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_545 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2301__A _2301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_589 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_56 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4334__CLK _4334_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4228__A _4247_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3132__A _3132_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_679 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2971__A _2953_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_44 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_392 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4484__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_554 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_205 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_227 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2756__A2 _2755_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_309 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_499 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_85 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_74 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3307__A _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2211__A _2210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_650 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_661 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3026__B _3105_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_397 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4130__A1 _4316_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_672 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2865__B _2865_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_624 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_698 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4138__A utmi_linestate_i[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3042__A _3041_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_167 VGND VPWR sky130_fd_sc_hd__fill_2
X_3920_ _3920_/A _2560_/X _3920_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_63_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_584 VGND VPWR sky130_fd_sc_hd__fill_2
X_3851_ _4534_/Q _3844_/X _3851_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2995__A2 _2993_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2802_ _2626_/Y _2638_/Y _2802_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3782_ _3785_/A _3782_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_81_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_615 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4304__C _2815_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2733_ _2733_/A _2727_/X _4215_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_117_147 VGND VPWR sky130_fd_sc_hd__fill_2
X_2664_ _2691_/A _2670_/B _2663_/X _2664_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_4403_ _4403_/D _4403_/Q _2411_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2595_ _2595_/A _2743_/A _2596_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_554 VGND VPWR sky130_fd_sc_hd__fill_1
X_4334_ _3288_/Y _2930_/A _2493_/X _4334_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2759__C _4469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3217__A _3146_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4558__RESET_B _2226_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_565 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_4265_ _4265_/A _4263_/X _4265_/C _4265_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4357__CLK _4356_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4196_ _4194_/Y _4196_/B _4199_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_3216_ _3216_/A _3216_/B _3216_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_82_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4048__A _4048_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3147_ _3041_/X _3151_/D _3146_/X _3228_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_27_326 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3880__B1 _3879_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_443 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_359 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3887__A _4549_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_627 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_679 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_167 VGND VPWR sky130_fd_sc_hd__fill_2
X_3078_ _3014_/Y _3037_/X _3188_/D _3077_/X _3132_/A VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__2791__A _2691_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_498 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3102__D _4359_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_381 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3699__B1 _3683_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4230__B _4276_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_180 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2669__C _2691_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3163__A2 _2999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2990__B1_N _2989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4112__A1 _4109_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3871__B1 _3870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_432 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_87 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_137 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_329 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3012__D _3011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_351 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2206__A _2206_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3926__A1 _2552_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_128 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3037__A _3019_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3154__A2 _3080_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2380_ _2379_/A _2380_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_312 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2876__A _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_440 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4103__B2 _4102_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2595__B _2743_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4050_ _4050_/A _4050_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3001_ _2886_/X _2906_/X _2850_/X _3277_/A VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_37_624 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3862__B1 _3861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_134 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3203__C _3203_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_167 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4470__SET_B _2330_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3500__A _3516_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3903_ _3884_/A _3897_/X _3902_/X _3903_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3090__A1 _3035_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3834_ _4519_/Q _3830_/X _3834_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_60_693 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2761__D _2760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_373 VGND VPWR sky130_fd_sc_hd__decap_8
X_3765_ _3762_/Y _3764_/X _3765_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_3696_ _3671_/X _3695_/B _3695_/X _3696_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__3393__A2 _3394_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2716_ _4497_/Q _2716_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2647_ _4527_/Q _2647_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4392__RESET_B _2423_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_49 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_673 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_340 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4321__RESET_B _2508_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2578_ _3925_/A _2578_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_101_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_524 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2786__A _2620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_237 VGND VPWR sky130_fd_sc_hd__fill_2
X_4317_ _2833_/X _4317_/Q _2512_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_101_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_345 VGND VPWR sky130_fd_sc_hd__decap_4
X_4248_ _2696_/A _4265_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_19_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_624 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2656__A1 _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_443 VGND VPWR sky130_fd_sc_hd__fill_2
X_4179_ _4179_/A _4180_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_27_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_646 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_24 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_156 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_679 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_318 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2959__A2 _2918_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3410__A _4368_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2671__D _2671_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_423 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4522__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4409__RESET_B _2404_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_489 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2592__B1 _4127_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_701 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4598__D _4212_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_535 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2696__A _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_53 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4097__B1 _4096_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_590 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_101 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_134 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_635 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_178 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2862__C _4404_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3320__A _3653_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4135__B _4135_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4021__B1 _4015_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3550_ _2865_/C _3541_/B _3550_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4151__A _4143_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2501_ _2497_/A _2501_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_3481_ _4421_/Q _3478_/B _3481_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3990__A _3990_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2432_ _2425_/A _2434_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_44_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2886__A1 _4375_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2363_ _2362_/A _2363_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_343 VGND VPWR sky130_fd_sc_hd__decap_8
X_4102_ _3915_/Y _4108_/B _3915_/Y _4108_/B _4102_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_398 VGND VPWR sky130_fd_sc_hd__fill_2
X_2294_ _2288_/X _2294_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4033_ _4033_/A _4033_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3835__B1 _3834_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_72 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4029__C _4029_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_649 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_608 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4545__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3884__B _3877_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3817_ _2658_/Y _3803_/X _3816_/X _3817_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_20_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4070__A1_N _4012_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_242 VGND VPWR sky130_fd_sc_hd__decap_3
X_3748_ _3749_/A _3747_/Y _3748_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4061__A _4061_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4502__RESET_B _2292_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_48 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_3679_ _3679_/A _3702_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_121_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3118__A2 _3094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3405__A _3402_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_207 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_711 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4236__A _4236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4023__A1_N _3969_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2682__C _2666_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_254 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3140__A _3036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_287 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_55 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_28 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4003__B1 _3972_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3357__A2 _3351_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_347 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_407 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3109__A2 _3375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_81 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_9 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2857__C _3563_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3315__A _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4418__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3817__B1 _3816_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_432 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_443 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_593 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_571 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_424 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4146__A _4137_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_468 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4568__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3050__A _3049_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2981_ _4429_/Q _3298_/B _4429_/Q _3298_/B _2981_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_21_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_3602_ _3585_/X _3602_/B _3601_/X _3602_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3348__A2 _3347_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4582_ _4582_/D _4582_/Q _2197_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_3533_ _3545_/A _3533_/B _3533_/C _3533_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3209__B _3205_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_29 VGND VPWR sky130_fd_sc_hd__decap_3
X_3464_ _3464_/A _3437_/B _3467_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_278 VGND VPWR sky130_fd_sc_hd__fill_2
X_2415_ _2411_/A _2415_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_440 VGND VPWR sky130_fd_sc_hd__fill_2
X_3395_ _3386_/X _3398_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3225__A _3077_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_162 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_2346_ _2339_/A _2352_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_516 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_207 VGND VPWR sky130_fd_sc_hd__fill_2
X_2277_ _2277_/A _2277_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3879__B _3877_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4016_ utmi_data_out_o[6] _4016_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_65_582 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4056__A _4079_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3895__A utmi_data_in_i[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4233__B1 _4612_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_438 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3110__D _3382_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2795__B1 _2794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_7 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3339__A2 _3326_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2304__A _2306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_584 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_317 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3119__B _3115_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_226 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3135__A _3055_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_685 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_560 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_585 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4495__RESET_B _2301_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4116__D _4116_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4424__RESET_B _2386_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_601 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_685 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2214__A _2210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_689 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_204 VGND VPWR sky130_fd_sc_hd__fill_1
X_2200_ _2199_/A _2200_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3045__A _3044_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3180_ _3136_/X _3176_/X _3077_/X _3179_/Y _3180_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_79_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_195 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2884__A _2872_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_132 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4390__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_327 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_2964_ _2955_/Y _2957_/Y _2960_/Y _2963_/Y _2964_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_22_449 VGND VPWR sky130_fd_sc_hd__decap_8
X_2895_ _3634_/A _3643_/A _4384_/Q _2894_/Y _2895_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2529__B1 _4616_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_82 VGND VPWR sky130_fd_sc_hd__decap_8
X_4565_ _4565_/D _4565_/Q _2218_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_116_565 VGND VPWR sky130_fd_sc_hd__fill_2
X_3516_ _3516_/A _3516_/B _3517_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3741__A2 _3740_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_204 VGND VPWR sky130_fd_sc_hd__decap_4
X_4496_ _4496_/D _4496_/Q _2300_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3447_ _4429_/Q _3434_/B _3450_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_85_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_600 VGND VPWR sky130_fd_sc_hd__fill_2
X_3378_ _2907_/X _3374_/X _3352_/Y _2851_/X _3377_/X _3379_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
X_2329_ _2330_/A _2329_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_270 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_493 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3105__D _3105_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_508 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3402__B _3398_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_379 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_224 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_449 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2768__B1 _4242_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_409 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4221__A3 _4116_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2963__A1_N _4421_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_392 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3732__A2 _3669_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4447__SET_B _2358_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_50 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_587 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2688__B _2674_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_408 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_471 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_368 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3799__A2 _3785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2209__A _2252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4127__C _4127_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4605__RESET_B _2170_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_703 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_585 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_276 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4606__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ _2680_/A _2679_/X _2680_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2879__A _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_497 VGND VPWR sky130_fd_sc_hd__fill_2
X_4350_ _3233_/Y _4350_/Q _2474_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_98_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_3301_ _3240_/A _3317_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4281_ _4281_/A _4282_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_4_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_681 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_460 VGND VPWR sky130_fd_sc_hd__fill_2
X_3232_ _2907_/X _3229_/Y _3412_/A _3232_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3206__C _3031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_3163_ _3920_/A _2999_/X _3240_/A _3163_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__3503__A _3503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_655 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_625 VGND VPWR sky130_fd_sc_hd__decap_12
X_3094_ _3359_/A _3359_/B _3021_/X _3105_/D _3094_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_81_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_390 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3222__B _3208_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_574 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4346__RESET_B _2479_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_511 VGND VPWR sky130_fd_sc_hd__decap_8
X_3996_ _4116_/D _3993_/B _3996_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2947_ _4428_/Q _2946_/X _4428_/Q _2946_/X _2947_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__4053__B _4053_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_318 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3693__A1_N _2650_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2789__A _4508_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2878_ _2877_/X _2878_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4617_ _4296_/Y _2524_/C _2154_/X _4619_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3714__A2 _3671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_502 VGND VPWR sky130_fd_sc_hd__decap_12
X_4548_ _3903_/X _3884_/A _2237_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4479_ _3743_/X _3709_/B _2320_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_104_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_268 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_666 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3413__A _3413_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_508 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4228__B _4228_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3132__B _3129_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2971__B _2964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_691 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_78 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_544 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_235 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_401 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2699__A _2624_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3166__B1 _3061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_467 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3307__B _2943_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_600 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3026__C _3350_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_538 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_30 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2865__C _2865_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3323__A _3317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4130__A2 _3960_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_463 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_614 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4138__B utmi_linestate_i[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_433 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_669 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_198 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_563 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_574 VGND VPWR sky130_fd_sc_hd__decap_4
X_3850_ _4525_/Q _3841_/X _3849_/X _3850_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4154__A _4153_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_555 VGND VPWR sky130_fd_sc_hd__fill_2
X_3781_ _3781_/A _3785_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_2801_ _2801_/A _2803_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_74_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4304__D _2824_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2732_ _2713_/X _2733_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3993__A _4116_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2663_ _2680_/A _2662_/X _2663_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3157__B1 _3055_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2402__A _2399_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4402_ _3533_/Y _2862_/A _2412_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2594_ _4050_/A _2743_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4333_ _3284_/Y _2928_/A _2494_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_577 VGND VPWR sky130_fd_sc_hd__fill_2
X_4264_ _3399_/A _4264_/B _4265_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_59_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_538 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_527 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4598__RESET_B _2178_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3215_ _4349_/Q _3216_/A VGND VPWR sky130_fd_sc_hd__inv_8
Xclkbuf_4_14_0_clk_i clkbuf_3_7_0_clk_i/X clkbuf_5_29_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_67_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3233__A _3231_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_132 VGND VPWR sky130_fd_sc_hd__decap_4
X_4195_ _4194_/Y _4196_/B _4197_/B VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3880__A1 _4538_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4527__RESET_B _2263_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_474 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4048__B _4073_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3146_ _3145_/X _3146_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_82_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_496 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_647 VGND VPWR sky130_fd_sc_hd__fill_2
X_3077_ _3059_/Y _3205_/C _3074_/X _3076_/X _3077_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3887__B _3895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_533 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_37 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3979_ _3994_/B _3979_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_109_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_58 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_47 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3699__A1 _3683_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2312__A _2314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3699__B2 _3698_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_310 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_205 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_459 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_430 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4112__A2 _4111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_411 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_33 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_22 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_305 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3871__A1 _4534_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4451__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2982__A _2940_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_99 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_628 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_691 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_319 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_54 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_544 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_599 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_396 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3926__A2 _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2222__A _2217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3037__B _3026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_286 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_717 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2876__B _4379_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4566__SET_B _2216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3053__A _3007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4149__A _4153_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_463 VGND VPWR sky130_fd_sc_hd__fill_2
X_3000_ _4231_/C _3003_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4620__RESET_B _4309_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3862__A1 _4530_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_282 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_146 VGND VPWR sky130_fd_sc_hd__decap_6
X_3902_ utmi_data_in_i[4] _3904_/B _3902_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_44_190 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3090__A2 _3088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_330 VGND VPWR sky130_fd_sc_hd__fill_2
X_3833_ _4517_/Q _3827_/X _3832_/X _3833_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_60_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_363 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3378__B1 _2851_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3764_ _3669_/C _3763_/X _3669_/C _3763_/X _3764_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3695_ _3695_/A _3695_/B _3695_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2715_ _2711_/X _2714_/X _2715_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_479 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_107 VGND VPWR sky130_fd_sc_hd__decap_8
X_2646_ _2645_/X _2646_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4324__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3228__A _3228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_363 VGND VPWR sky130_fd_sc_hd__decap_3
X_2577_ _2554_/X _2577_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_114_685 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4474__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_536 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2786__B _2810_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4316_ _2848_/X _4316_/Q _2513_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_249 VGND VPWR sky130_fd_sc_hd__decap_12
X_4247_ _4247_/A _4250_/B _4246_/X _4247_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__4059__A _4561_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_208 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4361__RESET_B _2461_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4178_ _4186_/B _4178_/B _4179_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3898__A utmi_data_in_i[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_591 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2656__A2 _2633_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_617 VGND VPWR sky130_fd_sc_hd__fill_2
X_3129_ _3129_/A _3112_/X _3119_/X _3181_/A _3129_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_82_285 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2307__A _2306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3410__B _3394_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_672 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_171 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_558 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_457 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_20_0_clk_i_A clkbuf_5_21_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_479 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2592__A1 _2566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_713 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3138__A _3227_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2696__B _2696_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__RESET_B _2356_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_61 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4097__A1 _4093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_282 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_20 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3601__A outport_data_o[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_617 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_263 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_116 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3057__C1 _3056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2862__D _4407_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_64 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3320__B _3320_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2217__A _2238_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_672 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4021__B2 _4020_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4347__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4151__B _4151_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2500_ _2497_/A _2500_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3480_ _3483_/A _3478_/Y _3480_/C _4420_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_6_562 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3048__A _3047_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_591 VGND VPWR sky130_fd_sc_hd__fill_2
X_2431_ _2431_/A _2431_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4497__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2887__A _2905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_300 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2886__A2 _2884_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2362_ _2362_/A _2362_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_37_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_121 VGND VPWR sky130_fd_sc_hd__fill_2
X_2293_ _2288_/X _2293_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4101_ _4566_/Q _4007_/X _3957_/Y _3966_/Y _4108_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_110_165 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_517 VGND VPWR sky130_fd_sc_hd__fill_2
X_4032_ _4010_/X _4031_/B _4030_/X _4031_/Y _4034_/B VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3835__A1 _4518_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_591 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_293 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3511__A _3514_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_19 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_193 VGND VPWR sky130_fd_sc_hd__decap_12
X_3816_ _3816_/A _3805_/X _3816_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3747_ _3746_/X _3747_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4061__B _4059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_438 VGND VPWR sky130_fd_sc_hd__fill_2
X_3678_ _2639_/X _3678_/B _3677_/X _3678_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_2629_ _2628_/X _2629_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_121_419 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4542__RESET_B _2244_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_344 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3405__B _3405_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_666 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_591 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3421__A _3420_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_572 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_116 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3140__B _3095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_266 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_23 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_480 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4252__A _4242_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4003__A1 _4002_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4003__B2 _3981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4402__D _3533_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_609 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_554 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2500__A _2497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_587 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_482 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2857__D _2856_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_75 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3315__B _2991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_377 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_539 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3817__A1 _2658_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3331__A _4376_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_200 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_414 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4146__B _4146_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2980_ _3297_/A _2935_/X _2979_/Y _3298_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_15_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_609 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_491 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_631 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4162__A _4187_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_653 VGND VPWR sky130_fd_sc_hd__decap_12
X_3601_ outport_data_o[3] _3592_/B _3601_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3753__B1 _3720_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4581_ _4151_/X _4581_/Q _2198_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3532_ _3503_/A _3541_/B _3533_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3209__C _3208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_3463_ _3483_/A _3463_/B _3462_/X _3463_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_6_392 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3506__A _3506_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2410__A _2396_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2414_ _2411_/A _2414_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3394_ _4260_/A _3394_/B _3394_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3225__B _3221_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_664 VGND VPWR sky130_fd_sc_hd__fill_2
X_2345_ _2345_/A _2345_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_496 VGND VPWR sky130_fd_sc_hd__fill_2
X_2276_ _2277_/A _2276_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_185 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_550 VGND VPWR sky130_fd_sc_hd__fill_2
X_4015_ _4011_/Y _4014_/X _4011_/Y _4014_/X _4015_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4512__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3241__A _3241_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_594 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_458 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4233__B2 _3407_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_406 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_469 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3895__B _3895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_620 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_631 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2795__A1 _2624_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4072__A utmi_data_out_o[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_697 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3744__B1 _2645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3119__C _3117_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_235 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2320__A _2318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3416__A _3416_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_290 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3135__B _3098_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_557 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_485 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_474 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_314 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4247__A _4247_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3151__A _3046_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_447 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_620 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_664 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_635 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_675 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_697 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_657 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4464__RESET_B _2337_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_167 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_428 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_351 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2230__A _2228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_227 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4535__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_260 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_185 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_163 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2884__B _2875_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_667 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_550 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4157__A _4187_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_723 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3061__A _3060_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_520 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3996__A _4116_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_406 VGND VPWR sky130_fd_sc_hd__fill_2
X_2963_ _4421_/Q _3261_/B _4421_/Q _3261_/B _2963_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__2405__A _2408_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2894_ _2893_/Y _2871_/B _2853_/D _2878_/Y _2894_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__2529__A1 _4615_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_61 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_18 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_511 VGND VPWR sky130_fd_sc_hd__decap_8
X_4564_ _4564_/D _4564_/Q _2219_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3515_ _4414_/Q _3512_/B _3517_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_116_544 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_417 VGND VPWR sky130_fd_sc_hd__fill_2
X_4495_ _4495_/D _4495_/Q _2301_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3236__A _3366_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3446_ _3424_/X _3446_/B _3445_/X _3446_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_97_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_130 VGND VPWR sky130_fd_sc_hd__fill_2
X_3377_ _3375_/A _3369_/Y _3376_/Y _3377_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_2328_ _2330_/A _2328_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_282 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4067__A _4073_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2259_ _2258_/A _2259_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_572 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_542 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_428 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2315__A _2314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2768__B2 _4490_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_247 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3965__B1 _2611_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_472 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4408__CLK _4410_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_522 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_148 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2688__C _2642_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3146__A _3145_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4558__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_22 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2985__A _2947_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_561 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_659 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3799__A3 _4495_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_158 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4127__D _4126_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_383 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_597 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3956__B1 _2611_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_236 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2225__A _2228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_704 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2879__B _4379_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3300_ _3279_/A _3300_/B _3300_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4280_ _2516_/X _4276_/B _4280_/C _4280_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_3_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_258 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_450 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2895__A _3634_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3231_ _2916_/Y _3228_/X _3230_/X _3231_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XANTENNA__4133__B1 _3979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_192 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3206__D _3114_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_3162_ _3392_/A _3240_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3503__B _3513_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2695__B1 _2804_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_317 VGND VPWR sky130_fd_sc_hd__fill_2
X_3093_ _3068_/X _3227_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_81_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_704 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_715 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_597 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_203 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4386__RESET_B _2431_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_247 VGND VPWR sky130_fd_sc_hd__decap_12
X_3995_ _3993_/X _3994_/X _2602_/X _4557_/D VGND VPWR sky130_fd_sc_hd__o21a_4
X_2946_ _3293_/A _2933_/X _2945_/Y _2946_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_13_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_308 VGND VPWR sky130_fd_sc_hd__decap_3
X_2877_ _2876_/X _2877_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xclkbuf_4_10_0_clk_i clkbuf_3_5_0_clk_i/X clkbuf_5_21_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4616_ _4616_/D _4616_/Q _2155_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4547_ _3901_/X _4547_/Q _2239_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_374 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_514 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4500__D _4500_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_525 VGND VPWR sky130_fd_sc_hd__decap_8
X_4478_ _3738_/X _3675_/B _2321_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_104_569 VGND VPWR sky130_fd_sc_hd__decap_8
X_3429_ _3429_/A _3430_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_634 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2686__B1 _2666_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_656 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3413__B _3657_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_47 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_678 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3132__C _3202_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_715 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2971__C _2967_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_534 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_523 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_180 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_12 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3938__B1 _2581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4380__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4260__A _4260_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2699__B _2689_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_446 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3166__B2 _3110_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3166__A1 _3070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4410__D _4410_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_366 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_630 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3026__D _3359_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4115__B1 _3990_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_239 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3604__A outport_data_o[4] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2865__D _4411_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_453 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3323__B _3322_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_412 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_467 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_670 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_383 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_501 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4154__B _4151_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3780_ _3707_/A _3780_/B _3781_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_2800_ _2797_/Y _2799_/Y _2800_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_44_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_2731_ _2537_/X _2730_/D _2731_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3993__B _3993_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_105 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4170__A _4188_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4401_ _4401_/D _3582_/A _2413_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2662_ _2657_/X _2658_/Y _2653_/A _2661_/X _2662_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_67_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3157__A1 _3059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_501 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4320__D _4320_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2593_ _4595_/Q _2595_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_534 VGND VPWR sky130_fd_sc_hd__fill_2
X_4332_ _4332_/D _2926_/A _2495_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_5_62 VGND VPWR sky130_fd_sc_hd__decap_3
X_4263_ _4263_/A _4263_/B _4263_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3514__A _3514_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3214_ _3367_/A _3397_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_79_291 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3233__B _3232_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4194_ _4591_/Q _4194_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_94_250 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_604 VGND VPWR sky130_fd_sc_hd__decap_6
X_3145_ _3079_/X _3144_/X _3145_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_27_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_317 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3880__A2 _3869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_125 VGND VPWR sky130_fd_sc_hd__fill_2
X_3076_ _3036_/X _3044_/X _3176_/A _3076_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_54_158 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4290__C1 _4289_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_361 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_512 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_49 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2977__A1_N _4427_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4042__C1 _4041_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_589 VGND VPWR sky130_fd_sc_hd__fill_2
X_3978_ _3978_/A _4116_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2929_ _2928_/X _2948_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_108_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3699__A2 _3698_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_661 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_427 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3424__A _3660_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_572 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3871__A2 _3869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_272 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_158 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_489 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4255__A _4265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_331 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4405__D _3542_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2503__A _2496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_254 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3037__C _3085_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_141 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_504 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_152 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3334__A _3333_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4149__B _4147_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3862__A2 _3855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_445 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_618 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_286 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4165__A _4164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_372 VGND VPWR sky130_fd_sc_hd__fill_2
X_3901_ _4547_/Q _3897_/X _3900_/X _3901_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__2822__B1 _2624_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_394 VGND VPWR sky130_fd_sc_hd__decap_8
X_3832_ _4518_/Q _3830_/X _3832_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3378__A1 _2907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3378__B2 _3377_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3509__A _4412_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3763_ _2659_/X _2660_/X _2659_/X _2660_/X _3763_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3694_ _3687_/Y _3693_/X _3687_/Y _3693_/X _3695_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__2413__A _2411_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2714_ _2587_/Y _2713_/X _2714_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_582 VGND VPWR sky130_fd_sc_hd__decap_4
X_2645_ _4523_/Q _2645_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3228__B _3227_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_4315_ enable_i utmi_xcvrselect_o[0] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_331 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4619__CLK _4619_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2576_ _2572_/X _2575_/X _2576_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2786__C _2786_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3244__A _2849_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_196 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_559 VGND VPWR sky130_fd_sc_hd__fill_2
X_4246_ _4233_/X _4235_/X _4239_/X _4245_/X _4246_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4059__B _4058_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_250 VGND VPWR sky130_fd_sc_hd__fill_2
X_4177_ _4186_/B _4178_/B _4181_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3898__B _3895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_721 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_423 VGND VPWR sky130_fd_sc_hd__decap_4
X_3128_ _3123_/X _3124_/X _3125_/X _3128_/D _3181_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_27_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_681 VGND VPWR sky130_fd_sc_hd__fill_2
X_3059_ _3058_/X _3059_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4330__RESET_B _2498_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_459 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_504 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_353 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_364 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_36 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3419__A _3419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_47 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4572__SET_B _2208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2323__A _2318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_469 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2592__A2 _2576_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3138__B _3095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_480 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_664 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_5_24_0_clk_i_A clkbuf_5_25_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4235__A2_N _4368_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2696__C _2695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_559 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_689 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4489__RESET_B _2308_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2993__A _2920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4097__A2 _4095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4418__RESET_B _2393_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_294 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_10 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3601__B _3592_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_404 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3057__B1 _3052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_150 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_81 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_92 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3329__A _4397_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4151__C _4150_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2233__A _2236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_480 VGND VPWR sky130_fd_sc_hd__fill_1
X_2430_ _2431_/A _2430_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_574 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2887__B _2886_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_504 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3064__A _3038_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2361_ _2362_/A _2361_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_559 VGND VPWR sky130_fd_sc_hd__decap_12
X_2292_ _2288_/X _2292_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4100_ _3918_/Y _4022_/X _3918_/Y _4022_/X _4100_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_689 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_389 VGND VPWR sky130_fd_sc_hd__decap_8
X_4031_ _4010_/X _4031_/B _4031_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3999__A _4602_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3835__A2 _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3511__B _3509_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2408__A _2408_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_415 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_448 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_492 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_481 VGND VPWR sky130_fd_sc_hd__decap_8
X_3815_ _2674_/Y _3803_/X _3814_/X _3815_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_20_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_200 VGND VPWR sky130_fd_sc_hd__fill_2
X_3746_ _3671_/X _4474_/Q _3739_/Y _3745_/Y _3746_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3239__A _3397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3771__A1 _3727_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_390 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4441__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3677_ _3677_/A _3676_/X _3677_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2628_ _2694_/A _2624_/A _2628_/C _2628_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_102_601 VGND VPWR sky130_fd_sc_hd__fill_1
X_2559_ _4489_/Q _4488_/Q _2522_/X _2525_/X _2559_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_114_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_483 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4591__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_4229_ _4278_/C _4278_/D _2730_/X _4276_/B VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4582__RESET_B _2197_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3702__A _3702_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_177 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3287__B1 _2930_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_529 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_581 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4511__RESET_B _2282_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2318__A _2318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_595 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_297 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_161 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_695 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4252__B _4263_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_356 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4003__A2 _3994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_200 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3149__A _3073_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_43 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_566 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_326 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3278__B1 _2926_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__A _3612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_389 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3817__A2 _3803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_9 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3331__B _4375_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2228__A _2228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_297 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4146__C _4620_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_256 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_481 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4464__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4162__B _4158_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_183 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_194 VGND VPWR sky130_fd_sc_hd__decap_4
X_3600_ _2859_/A _3589_/X _3602_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4580_ _4147_/X _4144_/A _2199_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3059__A _3058_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3531_ _3544_/B _3541_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3753__A1 _3745_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_214 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2898__A _2896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3209__D _3179_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_3462_ _3522_/A _3462_/B _3462_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3506__B _3513_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2413_ _2411_/A _2413_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_109 VGND VPWR sky130_fd_sc_hd__decap_8
X_3393_ _3342_/B _3394_/B _3392_/X _3393_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_97_621 VGND VPWR sky130_fd_sc_hd__decap_8
X_2344_ _2345_/A _2344_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3225__C _3224_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_453 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_378 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_507 VGND VPWR sky130_fd_sc_hd__fill_2
X_2275_ _2277_/A _2275_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3522__A _3522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_540 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_242 VGND VPWR sky130_fd_sc_hd__fill_2
X_4014_ utmi_data_out_o[5] _4066_/A utmi_data_out_o[5] _4066_/A _4014_/X VGND VPWR
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_223 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_554 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_418 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2795__A2 _2654_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_643 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_654 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4072__B _4072_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4503__D _3817_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_175 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_676 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3744__A1 _2646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_575 VGND VPWR sky130_fd_sc_hd__fill_2
X_3729_ _3730_/A _3730_/B _3729_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3744__B2 _2674_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3119__D _3118_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_707 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_7 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2601__A _2601_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_109 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3416__B _4514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_676 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3432__A _3431_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_326 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4337__CLK _4334_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_529 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4247__B _4250_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3151__B _3008_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_543 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4487__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_89 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_267 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_245 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_459 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4263__A _4263_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_120 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4413__D _3514_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3607__A _3607_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_82 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_93 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2511__A _2159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_64 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4433__RESET_B _2375_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_291 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_131 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_112 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2884__C _2883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3342__A _2867_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_679 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4157__B _4153_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_595 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3996__B _3993_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2962_ _4329_/Q _2920_/B _2961_/Y _3261_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_97_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4173__A _4164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_440 VGND VPWR sky130_fd_sc_hd__fill_2
X_2893_ _2880_/A _2893_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4323__D _2845_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_473 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2529__A2 _4614_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_495 VGND VPWR sky130_fd_sc_hd__decap_4
X_4563_ _4042_/X _4563_/Q _2220_/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3514_ _3514_/A _3512_/Y _3514_/C _3514_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3517__A _3514_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2421__A _2419_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4494_ _3798_/X _4494_/Q _2302_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_691 VGND VPWR sky130_fd_sc_hd__decap_12
X_3445_ _3510_/A _3437_/B _3445_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3236__B _3235_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4476__SET_B _2323_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3376_ _3376_/A _3376_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2327_ _2330_/A _2327_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3252__A _3265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_315 VGND VPWR sky130_fd_sc_hd__fill_2
X_2258_ _2258_/A _2258_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3111__C1 _3110_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4067__B _4065_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_595 VGND VPWR sky130_fd_sc_hd__fill_2
X_2189_ _2188_/X _2189_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_25_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_204 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4083__A utmi_data_out_o[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_259 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3965__A1 _2572_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3965__B2 _3964_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_350 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_617 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_534 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3427__A _3426_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2331__A _2324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2688__D _2652_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_440 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2985__B _2978_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4258__A _4265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_315 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_294 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3162__A _3392_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4408__D _4408_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_702 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_126 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_66 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_392 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_565 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2506__A _2504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_204 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_240 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3956__A1 _2571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3956__B2 _4048_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2241__A _2241_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4502__CLK _4450_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3337__A _2850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4614__RESET_B _2157_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_537 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_559 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_248 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2895__B _3643_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3230_ _3229_/Y _2916_/Y _2850_/X _3230_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4133__A1 _2575_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2695__A1 _2694_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4168__A _4168_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3161_ _3161_/A _3920_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_121_592 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3892__B1 _3891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_443 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3072__A _3072_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4318__D _2835_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3092_ _3176_/A _3059_/Y _3112_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_90_660 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2416__A _2411_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_524 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_237 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_259 VGND VPWR sky130_fd_sc_hd__decap_12
X_3994_ _3994_/A _3994_/B _4557_/Q _3994_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_2945_ _2935_/X _2945_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_50_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_2876_ _2876_/A _4379_/Q _2876_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_4615_ _4280_/Y _4615_/Q _2156_/X _4619_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_320 VGND VPWR sky130_fd_sc_hd__fill_1
X_4546_ _3899_/X _4546_/Q _2240_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3247__A _2917_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2151__A _2381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4355__RESET_B _2469_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_4477_ _3732_/X _3669_/C _2322_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_89_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_3428_ _3498_/A _3428_/B _3429_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_89_259 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2686__A1 _2684_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3359_ _3359_/A _3359_/B _3347_/Y _3361_/B VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__4078__A utmi_data_out_o[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2686__B2 _2670_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_167 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_318 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2326__A _2330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2971__D _2970_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3938__A1 _2605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3938__B2 _3937_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4525__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_46 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4260__B _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_320 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2699__C _2698_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_414 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3166__A2 _3363_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_22 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2996__A _2996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_708 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4115__A1 _3990_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4115__B2 _4002_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_570 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3604__B _3592_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_624 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3874__B1 _3873_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_424 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3620__A _4378_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_543 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2236__A _2236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4021__A1_N _4015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_513 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_535 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4051__B1 _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_2730_ _3810_/A _4504_/Q _2729_/X _2730_/D _2730_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_8_230 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_117 VGND VPWR sky130_fd_sc_hd__fill_1
X_2661_ _2645_/X _2649_/Y _2659_/X _2660_/X _2661_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4170__B _4167_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4400_ _3581_/Y _4400_/Q _2414_/X _4407_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3067__A _4356_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3157__A2 _3094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4601__D _4222_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2592_ _2566_/X _2576_/Y _4127_/C _2592_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4331_ _4331_/D _4331_/Q _2497_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_557 VGND VPWR sky130_fd_sc_hd__fill_2
X_4262_ _4610_/Q _4263_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_5_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3514__B _3512_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_3213_ _2999_/X _3209_/X _3212_/Y _3213_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_67_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_123 VGND VPWR sky130_fd_sc_hd__decap_3
X_4193_ _4197_/A _4196_/B _4192_/Y _4590_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_94_240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_167 VGND VPWR sky130_fd_sc_hd__fill_2
X_3144_ _4358_/Q _3010_/X _3381_/A _3008_/X _3144_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_48_690 VGND VPWR sky130_fd_sc_hd__decap_12
X_3075_ _3070_/X _3176_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3530__A _2862_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2944__A2_N _2943_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_137 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4290__B1 _2718_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_502 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4548__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_332 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_354 VGND VPWR sky130_fd_sc_hd__fill_2
X_3977_ _2552_/X _3969_/Y _3976_/X utmi_data_out_o[7] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4042__B1 _4033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_579 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4536__RESET_B _2251_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2928_ _2928_/A _2968_/A _2928_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_50_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_117 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4511__D _4512_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2859_ _2859_/A _2859_/B _2859_/C _2860_/C VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_117_640 VGND VPWR sky130_fd_sc_hd__decap_3
X_4529_ _4529_/D _4529_/Q _2261_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_2_439 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3705__A _3705_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_345 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_8 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clk_i clkbuf_4_9_0_clk_i/A clkbuf_4_8_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_105_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3828__A1_N _3822_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3440__A outport_data_o[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_479 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4255__B _4252_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_343 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_568 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4271__A _4265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_590 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4421__D _4421_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_109 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_673 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_150 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3037__D _3036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3615__A _3612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_461 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_126 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_159 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3350__A _3347_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4165__B _4163_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3900_ utmi_data_in_i[3] _3904_/B _3900_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2822__B2 _2821_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2822__A1 _2691_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3831_ _4517_/Q _3830_/X _3831_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3762_ _3668_/X _3762_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3378__A2 _3374_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4181__A _4201_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3509__B _3512_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4331__D _4331_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_437 VGND VPWR sky130_fd_sc_hd__decap_4
X_3693_ _2650_/Y _3692_/X _2650_/Y _3692_/X _3693_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_2713_ _2712_/X _2713_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_2644_ _2643_/Y _4524_/Q _2653_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_2575_ _2575_/A _4437_/Q _2575_/C _2575_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4314_ enable_i utmi_termselect_o VGND VPWR sky130_fd_sc_hd__buf_2
XANTENNA__3525__A _3554_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_505 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2786__D _2785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3244__B _3244_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3838__B1 _3837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_326 VGND VPWR sky130_fd_sc_hd__decap_4
X_4245_ _4240_/X _4241_/X _4245_/C _4244_/X _4245_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_59_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_240 VGND VPWR sky130_fd_sc_hd__decap_4
X_4176_ _4176_/A _4186_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3127_ _3050_/X _3103_/X _3045_/X _3223_/B _3128_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3260__A _3268_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4370__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_243 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_427 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_38 VGND VPWR sky130_fd_sc_hd__fill_2
X_3058_ _3359_/A _3360_/A _3021_/X _3347_/B _3058_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2813__A1 _2694_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4506__D _4306_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_332 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_663 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_140 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4015__B1 _4011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4370__RESET_B _2450_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_685 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4091__A _4079_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_516 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2604__A _2604_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_437 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3419__B _3528_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3435__A outport_data_o[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_676 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3829__B1 utmi_rxactive_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_624 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_85 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_28_0_clk_i_A clkbuf_5_29_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2993__B _2992_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_251 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_722 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4266__A _4266_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_627 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3170__A _3219_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_287 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_107 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3057__A1 _3219_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4416__D _3523_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4458__RESET_B _2345_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_693 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_82 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4006__B1 _2602_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_60 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2514__A _4620_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3329__B _3566_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3345__A _3337_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_602 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2664__B1_N _2663_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2360_ _2339_/A _2362_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_313 VGND VPWR sky130_fd_sc_hd__fill_2
X_2291_ _2288_/X _2291_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2740__B1 _2730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_145 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4393__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_20 VGND VPWR sky130_fd_sc_hd__fill_2
X_4030_ _4029_/X _4030_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_189 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_86 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4176__A _4176_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3080__A _3079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3511__C _3511_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_671 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_619 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4326__D _3250_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_170 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_641 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_471 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_713 VGND VPWR sky130_fd_sc_hd__decap_12
X_3814_ _3814_/A _3805_/X _3814_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2424__A _2381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_212 VGND VPWR sky130_fd_sc_hd__fill_2
X_3745_ _4474_/Q _3745_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3239__B _3236_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3771__A2 _3770_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_380 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_407 VGND VPWR sky130_fd_sc_hd__decap_12
X_3676_ _3669_/X _3672_/X _3676_/C _3675_/X _3676_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_2627_ _2626_/Y _2694_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_2558_ _4352_/Q _2908_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_0_707 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_173 VGND VPWR sky130_fd_sc_hd__fill_2
X_2489_ _2496_/A _2495_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_679 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_379 VGND VPWR sky130_fd_sc_hd__fill_2
X_4228_ _4247_/A _4228_/B _4604_/D VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3702__B _3701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3287__A1 _3280_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3287__B2 _3277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_424 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_690 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_221 VGND VPWR sky130_fd_sc_hd__fill_2
X_4159_ _4143_/X _4157_/Y _4158_/X _4583_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_28_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_619 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4551__RESET_B _2234_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_630 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2798__B1 _2633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_471 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_674 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2334__A _2337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_379 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3149__B _3114_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_289 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2970__B1 _3491_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2775__A2_N _2773_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_523 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3165__A _3108_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_335 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_clk_i clkbuf_2_2_0_clk_i/X clkbuf_3_5_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_87_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_508 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3278__B2 _3277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__B _3610_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3278__A1 _3251_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2509__A _2504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_585 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3331__C _2893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_243 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_438 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_663 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4609__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_162 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2244__A _2241_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3738__C1 _3737_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_688 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_699 VGND VPWR sky130_fd_sc_hd__decap_3
X_3530_ _2862_/A _3543_/B _3533_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3753__A2 _3752_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2898__B _2897_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3461_ outport_data_o[6] _3522_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3075__A _3070_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2412_ _2411_/A _2412_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_302 VGND VPWR sky130_fd_sc_hd__decap_3
X_3392_ _3392_/A _3391_/Y _3392_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_42_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_410 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_633 VGND VPWR sky130_fd_sc_hd__fill_2
X_2343_ _2345_/A _2343_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3225__D _3202_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_154 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3803__A _3804_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_476 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3522__B _3516_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_688 VGND VPWR sky130_fd_sc_hd__fill_2
X_2274_ _2253_/A _2277_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_711 VGND VPWR sky130_fd_sc_hd__decap_12
X_4013_ utmi_data_out_o[1] _4012_/Y utmi_data_out_o[1] _4012_/Y _4066_/A VGND VPWR
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__2419__A _2419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_254 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4218__B1 _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_405 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_7_0_clk_i clkbuf_4_3_0_clk_i/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_37_298 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_482 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2154__A _2155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_493 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_132 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_543 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3744__A2 _4524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_187 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2952__B1 _2951_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_3728_ _3674_/D _3727_/X _3674_/D _3727_/X _3730_/B VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
X_3659_ _3426_/Y _3528_/B _3660_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_114_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_537 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3713__A _3713_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_176 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_36 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2329__A _2330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_42 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4247__C _4246_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4209__B1 _4212_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_243 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3151__C _3369_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_46 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_522 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_438 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_276 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_577 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_408 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4263__B _4263_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_279 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_633 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_615 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_626 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2999__A _3216_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_32 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3607__B _3589_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2943__B1 _2942_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_397 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3623__A _3612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_327 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2239__A _2241_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3342__B _3342_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4402__RESET_B _2412_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4431__CLK _4430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_202 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_544 VGND VPWR sky130_fd_sc_hd__decap_3
X_2961_ _2922_/B _2961_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4173__B _4163_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4604__D _4604_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4581__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_493 VGND VPWR sky130_fd_sc_hd__decap_8
X_2892_ _2877_/X _2872_/D _2872_/B _2867_/X _2874_/A _2892_/Y VGND VPWR sky130_fd_sc_hd__o32ai_4
XFILLER_8_41 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2702__A _2595_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4562_ _4562_/D _4562_/Q _2221_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__3517__B _3517_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3513_ _3513_/A _3513_/B _3514_/C VGND VPWR sky130_fd_sc_hd__and2_4
X_4493_ _3797_/X _4493_/Q _2304_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_3444_ outport_data_o[2] _3510_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_6_191 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3533__A _3545_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3375_ _3375_/A _3369_/Y _3376_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_2326_ _2330_/A _2326_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_102 VGND VPWR sky130_fd_sc_hd__fill_2
X_2257_ _2258_/A _2257_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_124 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_338 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3111__B1 _3108_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4067__C _4066_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_28 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_2188_ _2166_/X _2188_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_92_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_706 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_16 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4083__B _4082_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_419 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_279 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4514__D _3828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3965__A2 _3963_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_452 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3708__A _3708_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_502 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2612__A _2611_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_546 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3427__B _3427_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4111__A2_N _4110_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_452 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3443__A _4428_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2985__C _2981_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_68 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_251 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_240 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4258__B _4258_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4454__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_596 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4274__A _2516_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_216 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_241 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4424__D _4424_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_430 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__A2 _3954_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_452 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4482__SET_B _2316_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3618__A _3617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_93 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3169__B1 _3014_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2522__A _4486_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_489 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3337__B _3336_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_673 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_590 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2895__C _4384_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3353__A _2867_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4133__A2 _4127_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_571 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_clk_i clkbuf_2_3_0_clk_i/A clkbuf_2_2_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_3160_ _3137_/X _3141_/X _3216_/B _3160_/D _3160_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3892__A1 _4543_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_496 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2695__A2 _3717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_658 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_647 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_3091_ _3148_/A _3208_/A _3089_/X _3091_/D _3129_/A VGND VPWR sky130_fd_sc_hd__or4_4
Xclkbuf_5_31_0_clk_i clkbuf_5_30_0_clk_i/A _4331_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_82_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_127 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_341 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4184__A _4201_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4334__D _3288_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3993_ _4116_/C _3993_/B _3993_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2944_ _3455_/A _2943_/X _3455_/A _2943_/X _2944_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__3528__A _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2875_ _2861_/X _2867_/X _2874_/Y _2875_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4204__A1_N _2718_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4327__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2432__A _2425_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4614_ _4614_/D _4614_/Q _2157_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_30_293 VGND VPWR sky130_fd_sc_hd__decap_8
X_4545_ _3896_/X _4545_/Q _2241_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3247__B _3266_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_4476_ _4476_/D _3668_/A _2323_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__4477__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_205 VGND VPWR sky130_fd_sc_hd__fill_2
X_3427_ _3426_/Y _3427_/B _3428_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4395__RESET_B _2420_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_102 VGND VPWR sky130_fd_sc_hd__decap_4
X_3358_ _3334_/X _3354_/X _2907_/X _3358_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__4324__RESET_B _2505_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_16 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4078__B _4076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_293 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_433 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2686__A2 _3713_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2309_ _2306_/A _2309_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4509__D _2665_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_455 VGND VPWR sky130_fd_sc_hd__fill_2
X_3289_ _3289_/A _3275_/B _3289_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_146 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_628 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_500 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4094__A _3966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_672 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_clk_i clkbuf_4_5_0_clk_i/A clkbuf_5_9_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_110_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_396 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_558 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_25 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3938__A2 _3935_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_36 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2342__A _2345_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3438__A _3424_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2699__D _2679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_343 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2996__B _2908_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_335 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4269__A _4237_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4115__A2 _4603_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_676 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3874__A1 _4535_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4419__D _3477_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_488 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_680 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3620__B _3620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2517__A _2516_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_683 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_599 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_81 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4051__A1 _4561_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4051__B2 _3964_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_619 VGND VPWR sky130_fd_sc_hd__decap_4
X_2660_ _2647_/Y _2660_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2252__A _2252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_264 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3067__B _3016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2591_ _2591_/A _2577_/Y utmi_txvalid_o _4127_/C VGND VPWR sky130_fd_sc_hd__nand3_4
X_4330_ _4330_/D _4330_/Q _2498_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_5_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_709 VGND VPWR sky130_fd_sc_hd__decap_4
X_4261_ _4265_/A _4261_/B _4261_/C _4609_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4179__A _4179_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3514__C _3514_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_508 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_208 VGND VPWR sky130_fd_sc_hd__decap_6
X_3212_ _3210_/Y _2999_/X _3412_/A _3212_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__3083__A _3082_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4329__D _4329_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_720 VGND VPWR sky130_fd_sc_hd__decap_4
X_4192_ _4185_/Y _4192_/B _4192_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_67_455 VGND VPWR sky130_fd_sc_hd__fill_2
X_3143_ _3029_/X _3061_/X _3142_/X _3143_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3078__C1 _3077_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3074_ _3068_/X _3070_/X _3065_/X _3073_/Y _3074_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3530__B _3543_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_447 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2427__A _2431_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_672 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4290__A1 _2548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_385 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3976_ _2579_/X _3976_/B _3976_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4042__A1 _4563_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2927_ _2926_/X _2968_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_388 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3258__A _4328_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2162__A _2163_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2858_ _3607_/A _2858_/B _4393_/Q _4392_/Q _2859_/C VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_116_140 VGND VPWR sky130_fd_sc_hd__fill_2
X_2789_ _4508_/Q _2790_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_116_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_4528_ _3857_/X _3837_/A _2262_/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4505__RESET_B _2289_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3705__B _3705_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4459_ _4521_/Q outport_data_o[1] _2344_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4089__A utmi_data_out_o[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_591 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_433 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_596 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_488 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_127 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2337__A _2337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_458 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_31 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4255__C _4254_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_97 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4271__B _4271_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3168__A _3219_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_162 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2800__A _2797_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3615__B _3613_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_316 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_241 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3631__A _3331_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_285 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2247__A _2248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_222 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3350__B _3347_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_661 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2822__A2 _2820_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_182 VGND VPWR sky130_fd_sc_hd__fill_2
X_3830_ _3824_/X _3830_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_60_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_3761_ _3726_/X _3715_/B _2687_/X _3760_/Y _3761_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3378__A3 _3352_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4181__B _4181_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4612__D _4271_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_2_0_clk_i_A clkbuf_5_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2712_ _4353_/Q _3417_/D _2712_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_9_562 VGND VPWR sky130_fd_sc_hd__fill_2
X_3692_ _3690_/A _3691_/A _3690_/Y _3730_/A _3692_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_72_3 VGND VPWR sky130_fd_sc_hd__decap_6
X_2643_ _4520_/Q _2643_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_114_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3806__A _3806_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2710__A _2539_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2574_ _2606_/C _2575_/C VGND VPWR sky130_fd_sc_hd__inv_8
X_4313_ _4313_/HI utmi_xcvrselect_o[1] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_114_633 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3525__B _3516_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_528 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3838__A1 _2673_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4244_ _4610_/Q _3399_/Y _4610_/Q _3399_/Y _4244_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_18 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3541__A _3513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_4175_ _4197_/A _4178_/B _4175_/C _4175_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__4515__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_274 VGND VPWR sky130_fd_sc_hd__fill_2
X_3126_ _3048_/Y _3150_/D _3223_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_639 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3260__B _3260_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_458 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_447 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2157__A _2155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_650 VGND VPWR sky130_fd_sc_hd__fill_2
X_3057_ _3219_/A _3045_/X _3052_/X _3056_/X _3188_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__2813__A2 _2633_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_480 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_694 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_182 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4082__A1_N _4018_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_697 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_163 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4091__B _4091_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4015__B2 _4014_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_539 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3774__B1 _3773_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4522__D _3843_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3959_ _3959_/A utmi_data_out_o[5] VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_109_416 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2620__A _4510_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_716 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_705 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_644 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4020__A1_N _4016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_614 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_259 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3829__A1 utmi_rxvalid_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_24 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_594 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3451__A _3451_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_425 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_639 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4266__B _4263_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_447 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3170__B _3122_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_469 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3057__A2 _3045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_428 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_491 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_83 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4282__A _4282_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_72 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4006__A1 _3993_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_50 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_174 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_clk_i clkbuf_2_0_0_clk_i/X clkbuf_4_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__4432__D _3463_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4498__RESET_B _2298_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3329__C _3329_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4427__RESET_B _2383_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_510 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_82 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3626__A _3612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2530__A _2522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3345__B _3344_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4538__CLK _4539_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2740__A1 _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_647 VGND VPWR sky130_fd_sc_hd__decap_3
X_2290_ _2288_/X _2290_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_1_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_701 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_263 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3361__A _2907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4607__D _4255_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_553 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_244 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_469 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_193 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4192__A _4185_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2705__A _2705_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3813_ _2646_/Y _3803_/X _3812_/X _3813_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_20_314 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4342__D _3239_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3744_ _2646_/Y _4524_/Q _2645_/X _2674_/Y _3749_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3756__B1 _4525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3239__C _3238_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_19 VGND VPWR sky130_fd_sc_hd__decap_4
X_3675_ _3709_/B _3675_/B _3713_/B _3711_/B _3675_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3536__A _3545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_419 VGND VPWR sky130_fd_sc_hd__decap_12
X_2626_ _4510_/Q _2626_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2440__A _2443_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_3_0_clk_i clkbuf_5_3_0_clk_i/A _4497_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_114_463 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_2557_ _2556_/X _2557_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_625 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_102 VGND VPWR sky130_fd_sc_hd__decap_8
X_2488_ _2485_/A _2488_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4227_ _2601_/X _4247_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3287__A2 _3285_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_723 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4517__D _3833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_4158_ _4187_/C _4153_/X _4158_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_11 VGND VPWR sky130_fd_sc_hd__decap_4
X_3109_ _3046_/X _3375_/A _3381_/A _3008_/X _3382_/A VGND VPWR sky130_fd_sc_hd__o22a_4
X_4089_ utmi_data_out_o[6] _4090_/B _4091_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_16_609 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_22 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_480 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2798__A1 _2694_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_247 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_15 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2615__A utmi_txvalid_o VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3995__B1 _2602_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_653 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_303 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4591__RESET_B _2186_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4520__RESET_B _2271_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2970__B2 _2969_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3446__A _3424_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2350__A _2352_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_41 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3165__B _3153_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_290 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_411 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4277__A _4615_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_488 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3278__A2 _3275_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__C _3611_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_561 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_200 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3181__A _3181_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_594 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_436 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_190 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4427__D _4427_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_564 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3331__D _3331_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_469 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2525__A _4487_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_269 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_93 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4608__RESET_B _2165_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_612 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3738__B1 _3719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_667 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_678 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2260__A _2253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4360__CLK _4334_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3356__A _3367_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3460_ _3460_/A _3437_/B _3463_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_6_395 VGND VPWR sky130_fd_sc_hd__fill_2
X_2411_ _2411_/A _2411_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3391_ _4257_/A _3394_/B _3391_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_2342_ _2345_/A _2342_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_35_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4187__A _4137_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2273_ _2272_/A _2273_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3091__A _3148_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4012_ utmi_data_out_o[2] _4012_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_5_10_0_clk_i_A clkbuf_4_5_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_361 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4337__D _3300_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_266 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4218__A1 _4281_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_597 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_247 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3977__B1 _3976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2435__A _2434_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4349__RESET_B _2476_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_533 VGND VPWR sky130_fd_sc_hd__fill_2
X_3727_ _3670_/Y _3679_/A _3705_/A _3702_/A _3727_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3136__A1_N _3041_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_588 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3266__A _4330_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2952__A1 _4330_/Q VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_26_0_clk_i clkbuf_4_13_0_clk_i/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__2170__A _2168_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_227 VGND VPWR sky130_fd_sc_hd__fill_1
X_3658_ _3244_/B _3657_/X _3585_/X _4374_/D VGND VPWR sky130_fd_sc_hd__o21a_4
X_3589_ _3610_/B _3589_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2609_ _2605_/X _2577_/Y _2608_/Y _4436_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3901__B1 _3900_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3713__B _3713_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_549 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_701 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_520 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_564 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_553 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_715 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4209__A1 _3984_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3151__D _3151_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2960__A1_N _4420_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_69 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2345__A _2345_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_589 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_612 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_450 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_483 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4383__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_605 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_188 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2943__A1 _3306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3176__A _3176_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_11 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_343 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3904__A utmi_data_in_i[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_645 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3623__B _3623_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_177 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_136 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_715 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_394 VGND VPWR sky130_fd_sc_hd__decap_3
X_2960_ _4420_/Q _3257_/B _4420_/Q _3257_/B _2960_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__2255__A _2258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4442__RESET_B _2364_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4173__C _4188_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2631__B1 _2804_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2891_ _2861_/X _2891_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_42_280 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_20 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_503 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4620__D _4620_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2702__B _4050_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4561_ _4561_/D _4561_/Q _2222_/X _4325_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__3086__A _3015_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3512_ _4413_/Q _3512_/B _3512_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3517__C _3517_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4492_ _4492_/D _4492_/Q _2305_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_569 VGND VPWR sky130_fd_sc_hd__decap_4
X_3443_ _4428_/Q _3434_/B _3446_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3814__A _3814_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3533__B _3533_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3374_ _3353_/Y _3342_/B _3374_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2325_ _2330_/A _2325_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_306 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_296 VGND VPWR sky130_fd_sc_hd__fill_2
X_2256_ _2258_/A _2256_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_497 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3111__A1 _3150_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_372 VGND VPWR sky130_fd_sc_hd__fill_2
X_2187_ _2183_/A _2187_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_25_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_180 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2774__A2_N _2766_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_394 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2165__A _2163_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2622__B1 _2669_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_420 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4530__D _4530_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2612__B _2554_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_528 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3724__A _3724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_14 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_clk_i clkbuf_4_1_0_clk_i/A clkbuf_5_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_115_580 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3443__B _3434_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2985__D _2984_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_335 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_604 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4258__C _4258_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_13 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_575 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4274__B _4272_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_545 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_353 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4063__C1 _4062_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_84 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_420 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2613__B1 _2612_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_239 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_413 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2803__A _2803_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3169__A1 _3021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3169__B2 _3051_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4440__D _2762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_652 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3634__A _3634_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2895__D _2894_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4233__A2_N _4257_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_475 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3892__A2 _3883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_486 VGND VPWR sky130_fd_sc_hd__fill_2
X_3090_ _3035_/X _3088_/Y _3085_/B _3091_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_81_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_383 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_320 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4184__B _4183_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_673 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4615__D _4280_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3992_ _2701_/A _3991_/X _4556_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_35_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_386 VGND VPWR sky130_fd_sc_hd__fill_2
X_2943_ _3306_/A _2940_/B _2942_/Y _2943_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_15_291 VGND VPWR sky130_fd_sc_hd__fill_2
X_2874_ _2874_/A _2874_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2713__A _2712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3528__B _3528_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4613_ _4274_/Y _4234_/A _2160_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_300 VGND VPWR sky130_fd_sc_hd__decap_6
X_4544_ _4544_/D _4544_/Q _2242_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4350__D _3233_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_366 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3544__A _3516_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4475_ _3718_/X _3667_/A _2325_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3426_ _3528_/D _3426_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_615 VGND VPWR sky130_fd_sc_hd__fill_1
X_3357_ _2851_/X _3351_/Y _3356_/X _3357_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__2686__A3 _2785_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2308_ _2306_/A _2308_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_626 VGND VPWR sky130_fd_sc_hd__fill_2
X_3288_ _3279_/A _3287_/Y _3288_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_2239_ _2241_/A _2239_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_681 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4364__RESET_B _2457_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3096__B1 _3095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_320 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2843__B1 _2842_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_394 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4094__B utmi_data_out_o[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_545 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4525__D _3850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_504 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3719__A _3704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3938__A3 _3936_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2623__A _4516_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3438__B _3434_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_405 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4421__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3454__A _3424_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2996__C _2995_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_399 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4269__B _4253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_655 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3874__A2 _3869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_125 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4571__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4285__A _4502_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_139 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_523 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4435__D _4435_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3629__A _3612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_711 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4051__A2 _3964_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_clk_i_A clkbuf_4_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_559 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2533__A _2532_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3067__C _3071_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_298 VGND VPWR sky130_fd_sc_hd__decap_8
X_2590_ _2589_/X utmi_txvalid_o VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3364__A _3039_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_4260_ _4260_/A _4264_/B _4261_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_4_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_250 VGND VPWR sky130_fd_sc_hd__fill_2
X_3211_ _3392_/A _3412_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4191_ _4185_/Y _4192_/B _4196_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_79_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_3142_ _3082_/X _3151_/D _3142_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_445 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_478 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2708__A _4503_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3078__B1 _3188_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4195__A _4194_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3073_ _3110_/C _3073_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_82_459 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4561__SET_B _2222_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4290__A2 _2718_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_353 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4110__A2_N _4562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4345__D _4345_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_301 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_19 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3539__A _3545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_345 VGND VPWR sky130_fd_sc_hd__decap_3
X_3975_ _2572_/X _3973_/Y _2611_/X _3974_/Y _3976_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__4042__A2 _4037_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2926_ _2926_/A _2965_/A _2926_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2443__A _2443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3258__B _3266_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2857_ _2857_/A _3559_/A _3563_/A _2856_/X _2857_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4444__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_2788_ _2788_/A _2796_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_686 VGND VPWR sky130_fd_sc_hd__fill_2
X_4527_ _3854_/X _4527_/Q _2263_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3274__A _3246_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4458_ _4520_/Q outport_data_o[0] _2345_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4594__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4089__B _4090_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_358 VGND VPWR sky130_fd_sc_hd__fill_2
X_3409_ _3406_/Y _3409_/B _3409_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4545__RESET_B _2241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_33 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_581 VGND VPWR sky130_fd_sc_hd__fill_2
X_4389_ _3602_/X _2859_/A _2428_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_607 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2618__A _4514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_692 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_651 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_684 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3449__A _3513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_356 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2353__A _2339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4271__C _4271_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3168__B _3036_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_581 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_653 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_642 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2800__B _2799_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3184__A _3181_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_697 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3615__C _3615_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3912__A _4553_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_467 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_456 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3631__B _3620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_404 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2528__A _2527_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_489 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4317__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_297 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3350__C _3350_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_665 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4467__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_334 VGND VPWR sky130_fd_sc_hd__fill_2
X_3760_ _3708_/A _3760_/B _3759_/Y _3760_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__2263__A _2261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_676 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3232__B1 _3412_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3359__A _3359_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_507 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_80 VGND VPWR sky130_fd_sc_hd__decap_4
X_2711_ _2710_/X _2711_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4181__C _4180_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_541 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_581 VGND VPWR sky130_fd_sc_hd__decap_4
X_3691_ _3691_/A _3730_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2642_ _2641_/Y _4525_/Q _2642_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_65_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_6_0_clk_i_A clkbuf_4_3_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_601 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3806__B _3805_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2710__B _2730_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2573_ _2555_/A _2575_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3094__A _3359_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4312_ _4312_/HI utmi_op_mode_o[1] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_99_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_4243_ _4242_/Y _3388_/A _4236_/Y _4260_/A _4245_/C VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3822__A _3822_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_306 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3838__A2 _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3299__B1 _3297_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4174_ _4188_/D _4169_/X _4175_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3541__B _3541_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_562 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_702 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2438__A _2434_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3125_ _3019_/Y _3026_/X _3095_/X _3125_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_67_297 VGND VPWR sky130_fd_sc_hd__decap_8
X_3056_ _3085_/A _3026_/X _3055_/X _3056_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_82_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_640 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3269__A _3265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2173__A _2168_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3774__A1 _3769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_39 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4091__C _4090_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3958_ _2578_/X _3956_/X _2552_/X _3957_/Y _3959_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_109_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3889_ _3889_/A _3895_/B _3889_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2909_ _2909_/A _3319_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2901__A _4427_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2620__B _2620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3829__A2 _3822_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_199 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3451__B _3434_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_264 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2348__A _2352_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_383 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_372 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_234 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4239__C1 _4238_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_651 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_470 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_654 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4282__B _4282_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4006__A2 _4005_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_40 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_676 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_367 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3329__D _2855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_595 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3626__B _3626_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4467__RESET_B _2334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2530__B _2525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_483 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3642__A _3662_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2740__A2 _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2258__A _2258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_562 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3361__B _3361_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_99 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_565 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_429 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_481 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_665 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4192__B _4192_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2705__B _2705_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_3812_ _3812_/A _3805_/X _3812_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_698 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_142 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3756__A1 _2658_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_326 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_3743_ _3726_/X _3709_/B _3719_/X _3742_/X _3743_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3756__B2 _2650_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_247 VGND VPWR sky130_fd_sc_hd__decap_12
X_3674_ _3715_/B _3674_/B _3674_/C _3674_/D _3676_/C VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__2721__A _2720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_269 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3536__B _3534_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2625_ _4449_/Q _2691_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_431 VGND VPWR sky130_fd_sc_hd__fill_2
X_2556_ _4489_/Q _4488_/Q _4486_/Q _2523_/Y _2556_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3552__A _3555_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2487_ _2485_/A _2487_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_359 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_540 VGND VPWR sky130_fd_sc_hd__fill_2
X_4226_ _4207_/X _4225_/Y _4603_/Q _4207_/X _4603_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3287__A3 _3286_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_573 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2168__A _2168_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4157_ _4187_/C _4153_/X _4157_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__3692__B1 _3690_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_510 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_201 VGND VPWR sky130_fd_sc_hd__fill_2
X_3108_ _3044_/X _3065_/X _3108_/X VGND VPWR sky130_fd_sc_hd__and2_4
Xclkbuf_5_22_0_clk_i clkbuf_5_22_0_clk_i/A _4430_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_55_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_4088_ utmi_data_out_o[5] _4087_/X _4090_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_28_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_3039_ _4358_/Q _3039_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2798__A2 _2692_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_492 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3995__A1 _3993_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4533__D _3868_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_153 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_214 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3446__B _3446_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4560__RESET_B _2223_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_13 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3462__A _3522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_68 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3278__A3 _3276_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3181__B _3181_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_404 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2806__A _2638_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_289 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_470 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_643 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_676 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4443__D _2756_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_698 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_635 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3738__A1 _3726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4505__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3637__A _2853_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2541__A _4499_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3356__B _3355_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_330 VGND VPWR sky130_fd_sc_hd__fill_2
X_2410_ _2396_/A _2411_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_108_280 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_291 VGND VPWR sky130_fd_sc_hd__decap_12
X_3390_ _3353_/Y _3394_/B _3389_/X _3390_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_2341_ _2345_/A _2341_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4081__A1_N _3949_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2272_ _2272_/A _2272_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_307 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4618__D _4618_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4187__B _4146_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3091__B _3208_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4011_ utmi_data_out_o[3] _4011_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_28_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_189 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_521 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_510 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_554 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_705 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4218__A2 _2546_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_373 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_513 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_215 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2716__A _4497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_470 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_5_14_0_clk_i_A clkbuf_4_7_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_259 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3977__A1 _2552_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4353__D _2890_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_451 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_440 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_602 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3733__A2_N _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_635 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4389__RESET_B _2428_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3547__A _3547_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3726_ _3708_/A _3726_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2451__A _2449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3266__B _3266_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2952__A2 _2922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4318__RESET_B _2511_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_239 VGND VPWR sky130_fd_sc_hd__fill_1
X_3657_ _2763_/A _2763_/B _3656_/Y _3657_/D _3657_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_3588_ _3587_/X _3610_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_2608_ _2566_/X _2607_/Y _2608_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3901__A1 _4547_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2539_ _4500_/Q _3818_/A _3812_/A _4505_/Q _2539_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_0_528 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_668 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_657 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3282__A _3243_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4528__D _3857_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_11 VGND VPWR sky130_fd_sc_hd__fill_1
X_4209_ _3984_/A _2704_/A _4212_/C _4209_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_28_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4209__A2 _2704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2626__A _4510_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_502 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4305__B1_N _4304_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_237 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4528__CLK _4539_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_646 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_495 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_668 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2957__A2_N _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3457__A _3547_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_52 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2361__A _2362_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3176__B _3073_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2943__A2 _2940_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3904__B _3904_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4288__A _2760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_668 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3623__C _3623_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3192__A _2999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_627 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4438__D _2592_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_521 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3920__A _3920_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_256 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2536__A _4505_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3408__B1 _3412_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4173__D _4188_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4081__B1 _3949_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2631__B2 _2670_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2631__A1 _2601_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2890_ _2852_/Y _2887_/X _2996_/A _2890_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2271__A _2272_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3367__A _3367_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4560_ _4560_/D _4560_/Q _2223_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4411__RESET_B _2401_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3086__B _3360_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3511_ _3514_/A _3509_/Y _3511_/C _4412_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_4491_ _4491_/D _4491_/Q _2306_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_548 VGND VPWR sky130_fd_sc_hd__fill_2
X_3442_ _3424_/X _3439_/Y _3441_/X _4427_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3814__B _3805_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3373_ _2851_/X _3370_/X _3372_/X _3373_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__4198__A _4592_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3533__C _3533_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2324_ _2324_/A _2330_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_465 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3830__A _3824_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2255_ _2258_/A _2255_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4348__D _3213_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_543 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3111__A2 _3107_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2186_ _2183_/A _2186_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2446__A _2425_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_513 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_i_A clk_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_376 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_579 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2622__A1 _2796_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3277__A _3277_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_476 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_498 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2181__A _2166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_3709_ _3713_/A _3709_/B _3709_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_107_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_559 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3724__B _3722_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_721 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_627 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_682 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_321 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2356__A _2358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4274__C _4273_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_557 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4350__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_708 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4063__B1 _4050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_96 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_2_0_clk_i_A clkbuf_3_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_410 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2613__A1 _2552_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2803__B _2802_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3187__A _3045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_436 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3169__A2 _3035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_487 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_642 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3915__A _4561_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3634__B _3620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_424 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_413 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3650__A _4376_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_137 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2266__A _2261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_395 VGND VPWR sky130_fd_sc_hd__decap_3
X_3991_ _3990_/Y _3979_/X _3937_/Y _3981_/X _3991_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_23_719 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_2942_ _2986_/B _2942_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2873_ _2872_/X _2874_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3097__A _3031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_251 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3528__C _3528_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4612_ _4271_/Y _4612_/Q _2161_/X _4612_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_312 VGND VPWR sky130_fd_sc_hd__decap_8
X_4543_ _3892_/X _4543_/Q _2243_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3825__A _3824_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4109__A1 _4009_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4474_ _4474_/D _4474_/Q _2326_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__3544__B _3544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_518 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3868__B1 _3867_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3425_ _3528_/C _3498_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_540 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_605 VGND VPWR sky130_fd_sc_hd__fill_2
X_3356_ _3367_/A _3355_/Y _3356_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_595 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2974__A1_N _2902_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3287_ _3280_/X _3285_/X _3286_/X _2930_/A _3277_/X _3287_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_2307_ _2306_/A _2307_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_2238_ _2238_/A _2241_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3560__A _3583_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4373__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4293__B1 _4247_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3096__A1 _3227_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_310 VGND VPWR sky130_fd_sc_hd__decap_4
X_2169_ _2168_/A _2169_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2843__A1 _4322_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2176__A _2177_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_354 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_685 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2904__A _2901_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_538 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4333__RESET_B _2494_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4541__D _3888_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3438__C _3437_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_428 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3735__A _3736_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_304 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_47 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3454__B _3451_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_623 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_634 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_435 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3470__A _3486_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_608 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_416 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4285__B _3816_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4284__B1 _2548_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_340 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_630 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_505 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_376 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_61 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3629__B _3627_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4451__D _2671_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_244 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_6_0_clk_i_A clkbuf_4_7_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3067__D _4355_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3645__A _3662_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_505 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3364__B _3364_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_538 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4396__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3210_ _4348_/Q _3210_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4190_ _4620_/D _4202_/D _4192_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_3141_ _3138_/X _3188_/A _3141_/C _3128_/D _3141_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3074__A1_N _3068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_295 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_159 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_254 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4275__B1 _4614_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3072_ _3072_/A _3110_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3078__A1 _3014_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4195__B _4196_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_641 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_630 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_170 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4027__B1 _3957_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_516 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2724__A _2724_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3974_ _3974_/A _3974_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3539__B _3537_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2925_ _2924_/X _2965_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_2856_ _4397_/Q _3566_/A _2856_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4361__D _4361_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_593 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3555__A _3555_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2787_ _2786_/X _2788_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_676 VGND VPWR sky130_fd_sc_hd__fill_2
X_4526_ _3852_/X _4526_/Q _2264_/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_104_337 VGND VPWR sky130_fd_sc_hd__fill_2
X_4457_ _2796_/A _3416_/A _2347_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_49_28 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_348 VGND VPWR sky130_fd_sc_hd__decap_3
X_3408_ _3407_/Y _3386_/X _3412_/A _3409_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3710__C1 _3709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_12 VGND VPWR sky130_fd_sc_hd__decap_12
X_4388_ _3599_/X _2859_/B _2429_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_424 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_413 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3290__A _3243_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3339_ _2851_/X _3326_/X _3338_/X _3339_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_100_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_276 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_49 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2618__B _2784_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4585__RESET_B _2193_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4514__RESET_B _2278_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4536__D _3876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_365 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_66 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_482 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2634__A _4516_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_549 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3449__B _3462_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_560 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3465__A outport_data_o[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_236 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_17_0_clk_i clkbuf_4_8_0_clk_i/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3184__B _3183_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_442 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_276 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2528__B _2525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_479 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_619 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_438 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4446__D _4446_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3350__D _3325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_600 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_376 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4009__B1 _4563_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_302 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_324 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3768__C1 _3767_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3232__A1 _2907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3359__B _3359_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2710_ _2539_/X _2730_/D _2710_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3690_ _3690_/A _3690_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2641_ _4521_/Q _2641_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3375__A _3375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2572_ _2571_/X _2572_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4311_ _4311_/HI utmi_dppulldown_o VGND VPWR sky130_fd_sc_hd__conb_1
XANTENNA__3094__B _3359_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_4242_ _4242_/A _4242_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_4_280 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_722 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3299__A1 _3280_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3299__B2 _3277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_210 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2719__A _2719_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4173_ _4164_/Y _4163_/C _4188_/C _4188_/D _4178_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_95_585 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_254 VGND VPWR sky130_fd_sc_hd__decap_12
X_3124_ _3227_/D _3080_/Y _3014_/Y _3124_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_48_490 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4356__D _3357_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_118 VGND VPWR sky130_fd_sc_hd__decap_4
X_3055_ _3054_/X _3055_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4411__CLK _4410_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_419 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_460 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_611 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_685 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2454__A _2456_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_357 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3269__B _2966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_3957_ _4566_/Q _3957_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_11_508 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3774__A2 _3772_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2908_ _2886_/X _2906_/X _2908_/C _2907_/X _2908_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_3888_ _4541_/Q _3883_/X _3887_/X _3888_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4561__CLK _4325_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3285__A _2930_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2901__B _4428_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2839_ _4320_/Q _2831_/X _2838_/X _4320_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_117_451 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_101 VGND VPWR sky130_fd_sc_hd__fill_2
X_4509_ _2665_/X _2818_/A _2284_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2734__B1 _2731_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2629__A _2628_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_276 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4239__B1 _4249_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_438 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_408 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_482 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4282__C _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_74 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2364__A _2362_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2973__B1 _2972_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_563 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_585 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3626__C _3625_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2530__C _2530_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_508 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3923__A _4570_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3642__B _3642_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_8 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2539__A _4500_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_12 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4436__RESET_B _2371_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_500 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3361__C _3361_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_70 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4434__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2274__A _2253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_633 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4584__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_132 VGND VPWR sky130_fd_sc_hd__fill_2
X_3811_ _2649_/Y _3803_/X _3810_/X _4500_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_176 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_204 VGND VPWR sky130_fd_sc_hd__decap_8
X_3742_ _3680_/Y _3740_/X _3741_/Y _3742_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3756__A2 _2659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_3673_ _3673_/A _3674_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_259 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3536__C _3536_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2624_ _2624_/A _3717_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_410 VGND VPWR sky130_fd_sc_hd__decap_8
X_2555_ _2555_/A _4437_/Q _2568_/B VGND VPWR sky130_fd_sc_hd__nand2_4
X_2486_ _2485_/A _2486_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_498 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3552__B _3550_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2449__A _2449_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4225_ _4224_/Y _4216_/B _4214_/Y _2745_/Y _4219_/D _4225_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_56_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_4156_ _4156_/A _4187_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_110_693 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3692__B2 _3730_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3692__A1 _3690_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_522 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_213 VGND VPWR sky130_fd_sc_hd__fill_2
X_3107_ _3068_/X _3151_/D _3107_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_28_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_408 VGND VPWR sky130_fd_sc_hd__fill_2
X_4087_ _3957_/Y _4007_/X _3957_/Y _4007_/X _4087_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_419 VGND VPWR sky130_fd_sc_hd__fill_2
X_3038_ _4360_/Q _3038_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_102_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_68 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2652__C1 _2651_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2184__A _2183_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3995__A2 _3994_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_441 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_132 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2912__A _2912_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_237 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_226 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2955__B1 _2954_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3446__C _3445_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_432 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3380__B1 _3337_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_58 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4457__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3462__B _3462_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2359__A _2358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_468 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3181__C _3216_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_682 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_235 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_449 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2806__B _2679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_121 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_482 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_485 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_198 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3918__A _4562_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3738__A2 _3675_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3637__B _3620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2946__B1 _2945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_353 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_386 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3653__A _3653_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4617__RESET_B _2154_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_413 VGND VPWR sky130_fd_sc_hd__fill_2
X_2340_ _2345_/A _2340_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_316 VGND VPWR sky130_fd_sc_hd__fill_2
X_2271_ _2272_/A _2271_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2269__A _2272_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_457 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3123__B1 _3150_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4187__C _4187_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4010_ _4008_/X _4009_/X _4008_/X _4009_/X _4010_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3091__C _3089_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_224 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_330 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2882__C1 _2879_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_544 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_558 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3977__A2 _3969_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_569 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_18_0_clk_i_A clkbuf_4_9_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2732__A _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_658 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3547__B _3544_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3725_ _3708_/X _3668_/X _3719_/X _3724_/Y _4476_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_20_179 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_579 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_191 VGND VPWR sky130_fd_sc_hd__fill_2
X_3656_ _2763_/C _3419_/A _3656_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3563__A _3563_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3587_ _3586_/X _3587_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4358__RESET_B _2464_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2607_ _2605_/X _2562_/X _2606_/X _2607_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__3901__A2 _3897_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2538_ _4501_/Q _3812_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3282__B _2949_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2179__A _2177_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_39 VGND VPWR sky130_fd_sc_hd__fill_2
X_2469_ _2472_/A _2469_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4208_ _4207_/X _2721_/X _3978_/A _4207_/X _4208_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_360 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_34 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_490 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_341 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2907__A _2849_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4139_ _4138_/X _4201_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_363 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4471__SET_B _2329_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4544__D _4544_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_430 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_2_0_clk_i_A clkbuf_2_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_463 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__A _2641_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3457__B _3462_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_86 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3473__A _3503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4288__B _4287_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_135 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3192__B _3191_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_190 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_341 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2817__A _2818_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_393 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3920__B _2560_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_363 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3408__A1 _3407_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_599 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4454__D _2682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_227 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4081__B2 _4566_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_463 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2631__A2 _3717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_71 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3648__A _3547_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_293 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2552__A _2552_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_444 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3367__B _3367_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_477 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3510_ _3510_/A _3513_/B _3511_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_7_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_499 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3086__C _3071_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4490_ _3794_/X _4490_/Q _2307_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3441_ _3506_/A _3437_/B _3441_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4451__RESET_B _2354_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3383__A _3366_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3372_ _3337_/Y _3371_/X _3367_/A _3372_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_40_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2323_ _2318_/A _2323_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_287 VGND VPWR sky130_fd_sc_hd__fill_2
X_2254_ _2258_/A _2254_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_341 VGND VPWR sky130_fd_sc_hd__fill_2
X_2185_ _2183_/A _2185_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_93_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_503 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_599 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4364__D _4364_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_366 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2622__A2 _2620_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3558__A _3583_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_591 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2462__A _2460_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4539__RESET_B _2248_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3708_ _3708_/A _3708_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_107_538 VGND VPWR sky130_fd_sc_hd__fill_2
X_3639_ _3662_/A _3637_/X _3639_/C _3639_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3724__C _3723_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3293__A _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4539__D _3882_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_477 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2637__A _4447_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_650 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_48 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_706 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4063__A1 _4568_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_208 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_233 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2613__A2 _2566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_244 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3468__A _3498_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_41 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2372__A _2367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3187__B _3085_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_i_A clkbuf_3_7_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3169__A3 _3055_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4299__A _4489_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_632 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3326__B1 _3347_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_665 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_433 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4449__D _2664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_606 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3931__A _3931_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_585 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_71 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3650__B _3646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2547__A _2520_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_366 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_344 VGND VPWR sky130_fd_sc_hd__fill_2
X_3990_ _3990_/A _3990_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2941_ _2941_/A _2986_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_15_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2282__A _2283_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_2872_ _2876_/A _2872_/B _2869_/Y _2872_/D _2872_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_4611_ _4268_/Y _4240_/A _2162_/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3097__B _3347_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3528__D _3528_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4542_ _3890_/X _4542_/Q _2244_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4473_ _4473_/D _3695_/A _2327_/X _4473_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__4109__A2 _4108_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_379 VGND VPWR sky130_fd_sc_hd__fill_2
X_3424_ _3660_/A _3424_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4002__A _4603_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3868__A1 _4533_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4359__D _3373_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_552 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_703 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3841__A _3883_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3355_ _3352_/Y _3354_/X _3366_/A _3355_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__4518__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_563 VGND VPWR sky130_fd_sc_hd__fill_2
X_2306_ _2306_/A _2306_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3286_ _3243_/B _2973_/X _3286_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_58_639 VGND VPWR sky130_fd_sc_hd__fill_2
X_2237_ _2236_/A _2237_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_469 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2457__A _2456_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_108 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4293__A1 _4616_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3096__A2 _3094_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_514 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_480 VGND VPWR sky130_fd_sc_hd__fill_2
X_2168_ _2168_/A _2168_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2843__A2 _2831_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_13 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_528 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_68 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3288__A _3279_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2904__B _2902_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2192__A _2188_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4373__RESET_B _2447_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_33 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2920__A _4329_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_418 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3735__B _3734_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3454__C _3453_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3308__B1 _3306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_585 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_628 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_679 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_13_0_clk_i_A clkbuf_3_6_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2367__A _2339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_428 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4285__C _4506_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_661 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4284__A1 _2533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_503 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_352 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_13_0_clk_i clkbuf_4_6_0_clk_i/X _4460_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_44_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_396 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_539 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3795__B1 _2657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_230 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_591 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3629__C _3628_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_561 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_234 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_285 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_296 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2830__A _2846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3645__B _3643_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_371 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3661__A _3528_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3140_ _3036_/X _3095_/X _3141_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2277__A _2277_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4275__A1 _4497_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3071_ _3071_/A _4355_/Q _3023_/Y _4357_/Q _3072_/A VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3078__A2 _3037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_288 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_653 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_483 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_314 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4027__B2 _4026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3786__B1 _3785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_185 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_358 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2724__B _2544_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3973_ _2605_/X _3970_/Y _3971_/X _2581_/X _3972_/Y _3973_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XANTENNA__3539__C _3539_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2924_ _4331_/Q _2951_/A _2924_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_550 VGND VPWR sky130_fd_sc_hd__fill_2
X_2855_ _2855_/A _2855_/B _3582_/A _4400_/Q _2855_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_117_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_600 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3555__B _3553_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4525_ _3850_/X _4525_/Q _2265_/X _4534_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2786_ _2620_/B _2810_/B _2786_/C _2785_/X _2786_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_116_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_4456_ _2827_/X _2763_/A _2348_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4340__CLK _4430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4387_ _4387_/D _2857_/A _2430_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3407_ _4270_/A _3407_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3710__B1 _3704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_24 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3571__A _3555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_572 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_561 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_701 VGND VPWR sky130_fd_sc_hd__fill_1
X_3338_ _3334_/X _3337_/Y _3240_/A _3338_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_85_211 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4490__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3290__B _2976_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3269_ _3265_/A _2966_/X _3269_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_105_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_672 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2187__A _2183_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_300 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_642 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2915__A _3244_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_78 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_377 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4552__D _4552_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4554__RESET_B _2230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3777__B1 _3720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_572 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2650__A _4526_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3764__A1_N _3669_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_64 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_168 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3701__B1 _3681_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_308 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3481__A _4421_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_572 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_701 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_244 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2528__C _2528_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_620 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_171 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2825__A _2620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_653 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_642 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_333 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_355 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4009__A1 _3933_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4009__B2 _3949_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_314 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4462__D _4524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3768__B1 _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_689 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3232__A2 _3229_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_369 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3359__C _3347_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2640_ _2628_/C _3707_/A _2639_/X _2680_/A VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__3656__A _2763_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4363__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2560__A _2559_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_554 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3375__B _3369_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2571_ _2610_/A _2571_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_336 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2988__A1_N _3460_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4310_ _4310_/HI utmi_dmpulldown_o VGND VPWR sky130_fd_sc_hd__conb_1
XANTENNA__3940__B1 _2611_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3094__C _3021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_509 VGND VPWR sky130_fd_sc_hd__fill_2
X_4241_ _4242_/A _3388_/Y _4266_/A _4267_/A _4241_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3299__A2 _3297_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3391__A _4257_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_691 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_222 VGND VPWR sky130_fd_sc_hd__decap_4
X_4172_ _4587_/Q _4188_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_96_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_266 VGND VPWR sky130_fd_sc_hd__fill_2
X_3123_ _3019_/Y _3122_/Y _3150_/D _3123_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_82_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3054_ _3381_/A _3038_/Y _3011_/X _3010_/X _3054_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_82_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4372__D _4303_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_634 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_196 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_678 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_144 VGND VPWR sky130_fd_sc_hd__fill_1
X_3956_ _2571_/X _3954_/X _2611_/X _4048_/A _3956_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_2907_ _2849_/A _2907_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3887_ _4549_/Q _3895_/B _3887_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3566__A _3566_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2470__A _2472_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_391 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2901__C _4429_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3285__B _3275_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2838_ inport_data_i[3] inport_accept_o _2838_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2769_ _4240_/A _4266_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4508_ _4508_/D _4508_/Q _2285_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2734__B2 _4215_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2734__A1 _2727_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_229 VGND VPWR sky130_fd_sc_hd__decap_12
X_4439_ _4439_/D _3925_/A _2368_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_120_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_606 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_520 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_200 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4547__D _3901_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_352 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4239__A1 _4234_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_119 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_269 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3998__B1 _2602_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_631 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_37 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2645__A _4523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_20 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2772__A2_N _2770_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_42 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4386__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_97 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4282__D _2546_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3476__A _3506_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2380__A _2379_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2973__A1 _2930_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_41 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_568 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3922__B1 _2581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_306 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_680 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3642__C _3641_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_542 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2539__B _3818_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_295 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_24 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4457__D _2796_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_512 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_597 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_545 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_247 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_642 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4405__RESET_B _2408_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3344__B1_N _3343_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2555__A _2555_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_280 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_645 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_81 VGND VPWR sky130_fd_sc_hd__decap_6
X_3810_ _3810_/A _3805_/X _3810_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_3741_ _3680_/Y _3740_/X _3708_/A _3741_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_32_166 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3386__A _3385_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_3672_ _3670_/Y _3679_/A _3671_/X _4472_/Q _3672_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2290__A _2288_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_362 VGND VPWR sky130_fd_sc_hd__decap_4
X_2623_ _4516_/Q _2624_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_111 VGND VPWR sky130_fd_sc_hd__decap_3
X_2554_ _2553_/X _2554_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3913__B1 _2581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_590 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_2485_ _2485_/A _2485_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3552__C _3552_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_339 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_4224_ _2753_/X _4224_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_110_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_715 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4367__D _3409_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4155_ _4143_/X _4153_/X _4154_/Y _4582_/D VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3692__A2 _3691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_19 VGND VPWR sky130_fd_sc_hd__fill_2
X_3106_ _3105_/X _3151_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_83_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_236 VGND VPWR sky130_fd_sc_hd__decap_4
X_4086_ _3939_/A _4056_/X _4050_/X _4085_/Y _4086_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_83_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2465__A _2460_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3037_ _3019_/Y _3026_/X _3085_/A _3036_/X _3037_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2652__B1 _2648_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_623 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_144 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3296__A _3279_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3939_ _3939_/A _4043_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2955__B2 _4418_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_400 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3380__A1 _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_447 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_704 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3181__D _3180_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_556 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2375__A _2379_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_280 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_604 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_40 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2946__A1 _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_383 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3653__B _3646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4401__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_560 VGND VPWR sky130_fd_sc_hd__decap_12
X_2270_ _2272_/A _2270_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_637 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3123__A1 _3019_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4187__D _4187_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3091__D _3091_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4551__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_394 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2882__B1 _2880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2285__A _2283_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_409 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_514 VGND VPWR sky130_fd_sc_hd__decap_12
X_3724_ _3724_/A _3722_/Y _3723_/X _3724_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4005__A _3994_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3655_ _3660_/A _3653_/Y _3654_/X _3655_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_9_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3844__A _3824_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2606_ _2575_/A _4437_/Q _2606_/C _2606_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3563__B _3566_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3586_ _3498_/A _3528_/D _3498_/C _3528_/B _3586_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_114_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_2537_ _4500_/Q _3818_/A _4501_/Q _3820_/A _2537_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4567__SET_B _2215_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_103 VGND VPWR sky130_fd_sc_hd__fill_2
X_2468_ _2496_/A _2472_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4398__RESET_B _2416_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4207_ _2706_/A _4207_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2399_ _2399_/A _2399_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4327__RESET_B _2501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_692 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_670 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_534 VGND VPWR sky130_fd_sc_hd__fill_2
X_4138_ utmi_linestate_i[1] utmi_linestate_i[0] _4138_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_589 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2195__A _2166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_409 VGND VPWR sky130_fd_sc_hd__decap_3
X_4069_ _3933_/Y _4022_/X _3933_/Y _4022_/X _4069_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_28_258 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2923__A _2922_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_272 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_637 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__B _4525_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_619 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_43 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4560__D _4560_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4424__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_313 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3473__B _3479_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_263 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4288__C _2533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4574__CLK _4574_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_266 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_480 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_139 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_225 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_707 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_386 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3408__A2 _3386_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2616__B1 _2591_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_90 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_291 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3929__A _4555_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2631__A3 _2691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_486 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3648__B _3646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_592 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_456 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4470__D _4470_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_67 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_630 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_140 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3086__D _3105_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_539 VGND VPWR sky130_fd_sc_hd__decap_3
X_3440_ outport_data_o[1] _3506_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_701 VGND VPWR sky130_fd_sc_hd__fill_1
X_3371_ _3334_/X _3342_/X _3371_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3344__A1 _3340_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3383__B _3381_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_712 VGND VPWR sky130_fd_sc_hd__decap_12
X_2322_ _2318_/A _2322_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_233 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4491__RESET_B _2306_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_158 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_266 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4420__RESET_B _2391_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2253_ _2253_/A _2258_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_320 VGND VPWR sky130_fd_sc_hd__fill_2
X_2184_ _2183_/A _2184_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_93_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3839__A _4529_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2607__B1 _2606_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_412 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2743__A _2743_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4447__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_283 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4380__D _3629_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_322 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3574__A _3516_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3707_ _3707_/A _3708_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_108_13 VGND VPWR sky130_fd_sc_hd__fill_2
X_3638_ outport_data_o[5] _3625_/B _3639_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4597__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_509 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_46 VGND VPWR sky130_fd_sc_hd__decap_4
X_3569_ _4397_/Q _3566_/B _3571_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3293__B _3275_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4579__RESET_B _2200_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_79 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4508__RESET_B _2285_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_288 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2918__A _4328_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_662 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_364 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4555__D _4555_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_718 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_567 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_386 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_239 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3749__A _3749_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_367 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4063__A2 _4056_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_234 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3271__B1 _4331_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_223 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2653__A _2653_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_389 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_581 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_245 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_53 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_456 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3484__A _3660_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4299__B _4488_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3326__B2 _3325_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_331 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2547__B _2546_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2837__B1 _2836_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4465__D _4527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_515 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4015__A2_N _4014_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__A _3426_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_654 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_2940_ _3306_/A _2940_/B _2941_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2563__A utmi_txready_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_209 VGND VPWR sky130_fd_sc_hd__fill_1
X_2871_ _2880_/A _2871_/B _2872_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_231 VGND VPWR sky130_fd_sc_hd__fill_2
X_4610_ _4265_/Y _4610_/Q _2163_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3097__C _3359_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4541_ _3888_/X _4541_/Q _2246_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3394__A _4260_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_460 VGND VPWR sky130_fd_sc_hd__fill_2
X_4472_ _4472_/D _4472_/Q _2328_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3423_ _3414_/A _3660_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_520 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3868__A2 _3855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4601__RESET_B _2175_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_220 VGND VPWR sky130_fd_sc_hd__fill_2
X_3354_ _3353_/Y _2857_/A _3354_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3285_ _2930_/A _3275_/B _3285_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2305_ _2306_/A _2305_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_618 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_106 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2738__A _2518_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2236_ _2236_/A _2236_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2828__B1 _4316_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4375__D _3649_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4293__A2 _3657_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_504 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_386 VGND VPWR sky130_fd_sc_hd__decap_8
X_2167_ _2166_/X _2168_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_81_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_25 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3569__A _4397_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_164 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2473__A _2472_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_209 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3288__B _3287_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2904__C _2904_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_581 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_18 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_152 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2920__B _2920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_336 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3308__B2 _3248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3308__A1 _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4342__RESET_B _2484_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2648__A _4523_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_117 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_128 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_109 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4612__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4284__A2 _4283_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_610 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_665 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_559 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3479__A _3510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2383__A _2388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_30 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3795__A1 _2684_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3795__B2 _3792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_573 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_268 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3645__C _3644_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_71 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3661__B _3498_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2558__A _4352_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_128 VGND VPWR sky130_fd_sc_hd__fill_2
X_3070_ _3069_/X _3070_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_94_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_662 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4275__A2 _2761_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_150 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2293__A _2288_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_676 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3235__B1 _3244_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_529 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3786__A1 _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_592 VGND VPWR sky130_fd_sc_hd__fill_2
X_3972_ _4560_/Q _3972_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2923_ _2922_/X _2951_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_540 VGND VPWR sky130_fd_sc_hd__decap_4
X_2854_ _2854_/A _2872_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_2785_ _2804_/A _4447_/Q _2785_/C _4450_/Q _2785_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_117_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3555__C _3554_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4524_ _3848_/X _4524_/Q _2266_/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_144 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_133 VGND VPWR sky130_fd_sc_hd__decap_4
X_4455_ _2671_/A _2620_/B _2349_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4386_ _3593_/X _2867_/A _2431_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3406_ _3607_/A _3398_/B _3406_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3710__A1 _3708_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3571__B _3571_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3337_ _2850_/X _3336_/X _3337_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2468__A _2496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_383 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_512 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_437 VGND VPWR sky130_fd_sc_hd__decap_12
X_3268_ _3268_/A _3268_/B _4330_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_85_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_407 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_470 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_150 VGND VPWR sky130_fd_sc_hd__decap_3
X_3199_ _3087_/X _3144_/X _3199_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_2219_ _2217_/X _2219_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_121_35 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2915__B _3241_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_183 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_389 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3777__A1 _3698_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_44 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2931__A _2930_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_595 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4594__RESET_B _2183_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4523__RESET_B _2268_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_21 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3762__A _3668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_411 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3701__B2 _3700_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3481__B _3478_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2378__A _2379_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_415 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_131 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2825__B _2800_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4009__A2 _4565_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3768__A1 _3724_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3002__A _3277_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4508__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_381 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3937__A _4556_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_511 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3656__B _3419_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_566 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2955__A2_N _4418_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_588 VGND VPWR sky130_fd_sc_hd__fill_2
X_2570_ _2552_/X _2554_/X _2569_/X _4439_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_114_626 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3672__A _3670_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3940__A1 _2572_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3940__B2 _4043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3094__D _3105_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_114 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_359 VGND VPWR sky130_fd_sc_hd__fill_2
X_4240_ _4240_/A _4240_/B _4240_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_4_293 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2288__A _2253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3299__A3 _3298_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3391__B _3394_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4171_ _4197_/A _4169_/X _4170_/Y _4171_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_95_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_532 VGND VPWR sky130_fd_sc_hd__decap_4
X_3122_ _3363_/A _3122_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_83_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_278 VGND VPWR sky130_fd_sc_hd__fill_2
X_3053_ _3007_/X _3381_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_36_621 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_109 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_473 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_484 VGND VPWR sky130_fd_sc_hd__decap_4
X_3955_ _3955_/A _4048_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3847__A _4532_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2906_ _2899_/Y _2905_/X _2906_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2751__A _2711_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3886_ _3824_/X _3895_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3566__B _3566_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2901__D _3451_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2837_ _4319_/Q _2831_/X _2836_/X _2837_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_2768_ _4242_/A _4490_/Q _4242_/A _4490_/Q _2768_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_117_475 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_615 VGND VPWR sky130_fd_sc_hd__fill_2
X_2699_ _2624_/A _2689_/B _2698_/X _2679_/X _2699_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_4507_ _2683_/X _2801_/A _2286_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2734__A2 _2730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_648 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3582__A _3582_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4438_ _2592_/Y _2591_/A _2369_/X _4574_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_120_618 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_381 VGND VPWR sky130_fd_sc_hd__decap_12
X_4369_ _3660_/Y _3528_/D _2451_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_86_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2198__A _2199_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_554 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4239__A2 _4368_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_364 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2926__A _2926_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_481 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3998__A1 _3996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_49 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_440 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_10 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4563__D _4042_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_646 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_32 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_175 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_657 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_359 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2661__A _2645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3476__B _3479_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2973__A2 _2948_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_514 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_464 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3922__A1 _2604_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3922__B2 _3921_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3492__A _3522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_329 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3686__B1 _2676_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2539__C _3812_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_554 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2836__A inport_data_i[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_654 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4473__D _4473_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_579 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2555__B _4437_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_153 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4330__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_101 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3667__A _3667_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3740_ _3671_/X _3687_/A _3739_/Y _3687_/Y _3740_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__2571__A _2610_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4445__RESET_B _2361_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3671_ _3695_/A _3671_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4480__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2622_ _2796_/A _2620_/X _2669_/A _2671_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_63_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_396 VGND VPWR sky130_fd_sc_hd__fill_2
X_2553_ _4620_/D utmi_txready_i _2553_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3913__B2 _3912_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3913__A1 _2604_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_478 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_145 VGND VPWR sky130_fd_sc_hd__decap_4
X_2484_ _2485_/A _2484_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_629 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_128 VGND VPWR sky130_fd_sc_hd__fill_2
X_4223_ _2704_/A _2733_/A _2754_/Y _4602_/Q _2706_/A _4602_/D VGND VPWR sky130_fd_sc_hd__a32o_4
X_4154_ _4153_/B _4151_/B _4154_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_110_684 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_587 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2746__A _4219_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4085_ _4079_/A _4083_/Y _4085_/C _4085_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_3105_ _3015_/X _4357_/Q _4354_/Q _3105_/D _3105_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_3036_ _3031_/X _3035_/X _3036_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3763__A1_N _2659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4383__D _3639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2652__A1 _2646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_421 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__A _3547_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_498 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_318 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2481__A _2475_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3296__B _3295_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3938_ _2605_/X _3935_/Y _3936_/X _2581_/X _3937_/Y _3938_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_3869_ _3883_/A _3869_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3701__A1_N _3681_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3380__A2 _3374_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4201__A _4201_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4558__D _4558_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_532 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_418 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_535 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4353__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4093__B1 _4568_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_462 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3840__B1 _3839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_145 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2391__A _2391_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3487__A _3504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_627 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2946__A2 _2933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_362 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_209 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_261 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4468__D _2826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_572 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_448 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3123__A2 _3122_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_384 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2566__A _2565_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2882__A1 _2878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_440 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_443 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3397__A _3397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_537 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_526 VGND VPWR sky130_fd_sc_hd__fill_1
X_3723_ _3670_/Y _3723_/B _3723_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4005__B _4552_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_3654_ _3554_/A _3646_/Y _3654_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2605_ _2604_/X _2605_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3585_ _3415_/Y _3585_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2536_ _4505_/Q _3820_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_0_509 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_415 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_115 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4378__D _3623_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2771__A2_N _4494_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2467_ _2381_/A _2496_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2570__B1 _2569_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_297 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4376__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4206_ _4205_/X _4212_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_2398_ _2399_/A _2398_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_705 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_14 VGND VPWR sky130_fd_sc_hd__fill_2
X_4137_ _2628_/C _4137_/B _4137_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2476__A _2475_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_568 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4075__B1 _3941_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4068_ _4569_/Q _4056_/X _4050_/X _4067_/Y _4068_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_83_387 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_29 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4367__RESET_B _2454_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_229 VGND VPWR sky130_fd_sc_hd__decap_8
X_3019_ _3018_/X _3019_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_616 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3100__A _3227_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_22 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_671 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_220 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_223 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3770__A _3727_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_107 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_470 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2386__A _2388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_52 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_557 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_719 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2616__A1 utmi_txready_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_410 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3813__B1 _3812_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_240 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3010__A _3009_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4573__SET_B _2207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4106__A _4079_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_435 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3945__A _4347_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_620 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_507 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4399__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_163 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3344__A2 _3342_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3370_ _3369_/A _3369_/B _3369_/Y _3370_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3383__C _3383_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_2321_ _2318_/A _2321_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3680__A _4472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_608 VGND VPWR sky130_fd_sc_hd__fill_2
X_2252_ _2252_/A _2253_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_2_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_671 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2296__A _2324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_535 VGND VPWR sky130_fd_sc_hd__decap_6
X_2183_ _2183_/A _2183_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4057__B1 _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4460__RESET_B _2343_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_313 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_376 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2607__A1 _2605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_207 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3839__B _3830_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_590 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2743__B _4443_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4016__A utmi_data_out_o[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_424 VGND VPWR sky130_fd_sc_hd__decap_3
X_3706_ _3705_/A _3705_/B _3704_/X _3705_/Y _4470_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__3855__A _3883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3574__B _3583_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_25 VGND VPWR sky130_fd_sc_hd__fill_2
X_3637_ _2853_/D _3620_/B _3637_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_103_702 VGND VPWR sky130_fd_sc_hd__fill_2
X_3568_ _3555_/A _3566_/Y _3567_/X _3568_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_103_713 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_18 VGND VPWR sky130_fd_sc_hd__fill_2
X_2519_ _2518_/X _2519_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3499_ _3498_/X _3516_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3590__A _2867_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4548__RESET_B _2237_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_267 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2918__B _2918_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_619 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4296__B1 _4295_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_502 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_674 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2934__A _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3271__A1 _3251_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3271__B2 _3248_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_224 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3749__B _3747_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_202 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2653__B _2652_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_560 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4571__D _4571_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_235 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_722 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_424 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_435 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_479 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3765__A _3762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4220__B1 _3990_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4541__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_551 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4299__C _2527_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_446 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_449 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_129 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2837__A1 _4319_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_641 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3005__A _3005_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_387 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_72 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2844__A inport_data_i[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__B _3528_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_677 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4481__D _4481_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2870_ _3331_/D _2871_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_43_593 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_60 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__A _3709_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_93 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3097__D _3359_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_4540_ _4540_/D _4540_/Q _2247_/X _4545_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4471_ _4471_/D _3679_/A _2329_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_116_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3394__B _3394_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_472 VGND VPWR sky130_fd_sc_hd__fill_2
X_3422_ _4372_/Q _3415_/Y _3422_/C _3422_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_112_532 VGND VPWR sky130_fd_sc_hd__decap_8
X_3353_ _2867_/A _3353_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_254 VGND VPWR sky130_fd_sc_hd__fill_2
X_3284_ _3279_/A _3283_/Y _3284_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_2304_ _2306_/A _2304_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2738__B _2546_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2235_ _2236_/A _2235_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_449 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_438 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2828__A1 _2557_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2166_ _2252_/A _2166_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4414__CLK _4410_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_622 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_685 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_674 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_173 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_162 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_644 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_184 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3569__B _3566_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_176 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4391__D _3609_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_593 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4564__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3585__A _3415_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_287 VGND VPWR sky130_fd_sc_hd__decap_8
X_2999_ _3216_/B _2999_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_131 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2764__B1 _4234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_359 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_28 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3308__A2 _3306_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_521 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2929__A _2928_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_637 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2648__B _4527_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_449 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_438 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4382__RESET_B _2436_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4566__D _4049_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_408 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_65 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_527 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3479__B _3479_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_165 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_700 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3795__A2 _3782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_715 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3495__A _3554_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_596 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2755__B1 _2754_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_442 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3914__A2_N _3913_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_381 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_395 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4476__D _4476_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4437__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4275__A3 _3657_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_82 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2574__A _2606_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4587__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_143 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3235__A1 _3319_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3971_ _3229_/Y _4278_/C _3971_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_16_560 VGND VPWR sky130_fd_sc_hd__decap_4
X_2922_ _4330_/Q _2922_/B _2922_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3786__A2 _3790_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_571 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2994__B1 _2850_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_390 VGND VPWR sky130_fd_sc_hd__fill_2
X_2853_ _3634_/A _3643_/A _4384_/Q _2853_/D _2854_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_31_585 VGND VPWR sky130_fd_sc_hd__decap_6
X_2784_ _2784_/A _4449_/Q _2696_/B _2786_/C VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_116_101 VGND VPWR sky130_fd_sc_hd__decap_4
X_4523_ _3846_/X _4523_/Q _2268_/X _4539_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_104_318 VGND VPWR sky130_fd_sc_hd__fill_2
X_4454_ _2682_/X _2696_/B _2350_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4385_ _3645_/X _3643_/A _2433_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3405_ _3402_/Y _3405_/B _3405_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2749__A _4501_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3710__A2 _3679_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3571__C _3571_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_3336_ _2896_/A _4375_/Q _3335_/Y _3336_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_112_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_37 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_235 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4386__D _3593_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_449 VGND VPWR sky130_fd_sc_hd__decap_3
X_3267_ _3251_/X _3265_/X _3266_/X _4330_/Q _3248_/X _3268_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_105_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_663 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_162 VGND VPWR sky130_fd_sc_hd__fill_2
X_3198_ _3019_/Y _3107_/Y _3085_/B _3198_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_2218_ _2217_/X _2218_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_493 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2484__A _2485_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_688 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4076__A2_N _4075_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_485 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3777__A2 _3776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_112 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2737__B1 _2736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4014__A2_N _4066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_137 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_189 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4477__SET_B _2322_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2659__A _4526_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_235 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_408 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_600 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_151 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2394__A _2391_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_463 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2825__C _2825_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3768__A2 _3674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_669 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2976__B1 _2975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3953__A _4348_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3940__A2 _3938_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3672__B _3679_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_349 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_714 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_4170_ _4188_/C _4167_/B _4170_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_3121_ _3120_/X _3363_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_121_192 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_408 VGND VPWR sky130_fd_sc_hd__fill_2
X_3052_ _3048_/Y _3051_/Y _3052_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_48_482 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_452 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_441 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_282 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_260 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_124 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_338 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_349 VGND VPWR sky130_fd_sc_hd__fill_2
X_3954_ _2581_/A _3952_/X _3953_/X _2604_/X _4558_/Q _3954_/X VGND VPWR sky130_fd_sc_hd__o32a_4
X_3885_ _4540_/Q _3883_/X _3884_/X _4540_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3847__B _3844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2967__B1 _3488_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2905_ _2905_/A _4418_/Q _2900_/X _2904_/X _2905_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2751__B _2750_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2836_ inport_data_i[2] inport_accept_o _2836_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4024__A _4564_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_454 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_443 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_421 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3863__A _4539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2767_ _4612_/Q _2765_/Y _4608_/Q _2766_/Y _2767_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4602__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2698_ _2654_/X _2662_/X _2698_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4506_ _4306_/Y _4506_/Q _2287_/X _4450_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_498 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3582__B _3582_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2479__A _2475_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4437_ _2603_/X _4437_/Q _2370_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_25 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3696__B1_N _3695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_224 VGND VPWR sky130_fd_sc_hd__fill_2
X_4368_ _3412_/Y _4368_/Q _2452_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_86_544 VGND VPWR sky130_fd_sc_hd__decap_8
X_3319_ _3319_/A _3320_/B _3319_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4299_ _4489_/Q _4488_/Q _2527_/Y _2523_/Y _4299_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_100_387 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2926__B _2965_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3998__A2 _3997_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3103__A _3102_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_22 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_102 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_33 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_187 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_55 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2942__A _2986_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_88 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_146 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_77 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2661__B _2649_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_99 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_10 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_382 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_599 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_476 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3922__A2 _3919_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2389__A _2396_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3492__B _3486_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3686__A1 _2646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_360 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2539__D _4505_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_192 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2836__B inport_accept_o VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_633 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_441 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_603 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_677 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3013__A _3012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_474 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_72 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2852__A _4353_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2949__B1 _2948_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_477 VGND VPWR sky130_fd_sc_hd__fill_1
X_3670_ _3705_/A _3670_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3683__A _3683_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2621_ _2601_/A _2669_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4414__RESET_B _2398_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2552_ _2552_/A _2552_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3913__A2 _3910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_435 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2299__A _2301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_2483_ _2485_/A _2483_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4222_ _4116_/D _4207_/X _4222_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_68_500 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_490 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_544 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_533 VGND VPWR sky130_fd_sc_hd__fill_1
X_4153_ _4153_/A _4153_/B _4147_/C _4153_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_110_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2746__B _4469_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3104_ _3103_/X _3150_/D VGND VPWR sky130_fd_sc_hd__inv_8
X_4084_ utmi_data_out_o[5] _4082_/X _4085_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_83_547 VGND VPWR sky130_fd_sc_hd__fill_2
X_3035_ _3359_/A _3360_/A _3347_/B _3035_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_36_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3115__A2_N _3018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_591 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_580 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2652__A2 _2647_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_474 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3858__A _3824_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_455 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_433 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2762__A _2757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__B _3583_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3937_ _4556_/Q _3937_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_23_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_691 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_218 VGND VPWR sky130_fd_sc_hd__decap_8
X_3868_ _4533_/Q _3855_/X _3867_/X _3868_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_3799_ _2601_/X _3785_/X _4495_/Q _4525_/Q _3792_/A _4495_/D VGND VPWR sky130_fd_sc_hd__a32o_4
X_2819_ _2639_/X _2698_/X _2819_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3593__A _3585_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_13 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_35 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_529 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_457 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_28 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_8 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4201__B _4199_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_544 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2937__A _2936_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_599 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_385 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_227 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4574__D _4098_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4093__B2 utmi_data_out_o[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4093__A1 _3969_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3840__A1 _2657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2672__A _2785_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_647 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3487__B _3485_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_477 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_168 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_341 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_352 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_323 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_617 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3008__A _4360_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_7 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_205 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4484__D _3775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2882__A2 _2861_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_536 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_525 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_558 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_528 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3678__A _2639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2582__A _2581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_252 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3397__B _3394_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_639 VGND VPWR sky130_fd_sc_hd__fill_2
X_3722_ _3670_/Y _3723_/B _3722_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_3653_ _3653_/A _3646_/Y _3653_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4302__A enable_i VGND VPWR sky130_fd_sc_hd__diode_2
X_2604_ _2604_/A _2604_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3584_ _3581_/A _3582_/Y _3583_/X _4401_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_2535_ _4504_/Q _3818_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2570__A1 _2552_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_276 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_127 VGND VPWR sky130_fd_sc_hd__decap_8
X_2466_ _2460_/X _2466_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_149 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2757__A _2716_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4205_ _2706_/A _2754_/Y _4205_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_2397_ _2399_/A _2397_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_650 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_91 VGND VPWR sky130_fd_sc_hd__decap_4
X_4136_ _4135_/B _4137_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_28_205 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4394__D _3562_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3684__A2_N _3669_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_355 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_506 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4075__B2 _4565_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4067_ _4073_/A _4065_/Y _4066_/X _4067_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_83_399 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_720 VGND VPWR sky130_fd_sc_hd__decap_4
X_3018_ _3017_/X _3018_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3588__A _3587_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2492__A _2495_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_230 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_422 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4336__RESET_B _2491_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3100__B _3084_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_650 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3338__B1 _3240_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4212__A _4210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4569__D _4068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_359 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_287 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4320__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3770__B _3770_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2667__A _2785_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_661 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4470__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_344 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3813__A1 _2646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_219 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2616__A2 _4029_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_271 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3498__A _3498_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_52 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_252 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__B _4104_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_425 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_650 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3945__B _3417_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4122__A _2605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_687 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4479__D _3743_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3961__A _3216_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_2320_ _2318_/A _2320_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2251_ _2248_/A _2251_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_127 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2577__A _2554_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2182_ _2183_/A _2182_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_333 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4057__A1 _3974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3700__A1_N _3682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4057__B2 utmi_data_out_o[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_219 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2607__A2 _2562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_282 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3201__A _3209_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_302 VGND VPWR sky130_fd_sc_hd__decap_3
X_3705_ _3705_/A _3705_/B _3705_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_107_519 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4343__CLK _4325_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3636_ _3662_/A _3634_/X _3636_/C _3636_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_3567_ _3510_/A _3582_/B _3567_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4389__D _3602_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_563 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3740__B1 _3739_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_202 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_403 VGND VPWR sky130_fd_sc_hd__fill_2
X_2518_ _3416_/A _4514_/Q _2763_/A _2518_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_115_596 VGND VPWR sky130_fd_sc_hd__fill_2
X_3498_ _3498_/A _3498_/B _3498_/C _3498_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3590__B _3589_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4493__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2487__A _2485_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2449_ _2449_/A _2449_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_661 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4296__A1 _2725_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_4119_ _3993_/B _4118_/X _4119_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_29_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_325 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4588__RESET_B _2190_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_208 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4517__RESET_B _2275_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2934__B _2933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_720 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3271__A2 _3269_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_252 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4207__A _2706_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_66 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_447 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3765__B _3764_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4220__B2 _4207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4220__A1 _2704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_491 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4299__D _2523_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_414 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3781__A _3781_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_555 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2397__A _2399_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_439 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_480 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2837__A2 _2831_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_40 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2844__B _2846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_689 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3798__B1 _4524_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_550 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3021__A _3071_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_572 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2860__A _2855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4366__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__B _3675_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_83 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4470_ _4470_/D _3705_/A _2330_/X _4470_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3421_ _3420_/X _3422_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_500 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3691__A _3691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_712 VGND VPWR sky130_fd_sc_hd__decap_12
X_3352_ _3334_/X _3352_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2303_ _2324_/A _2306_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_690 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_406 VGND VPWR sky130_fd_sc_hd__decap_4
X_3283_ _3280_/X _3281_/X _3282_/X _2928_/A _3277_/X _3283_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_58_609 VGND VPWR sky130_fd_sc_hd__decap_6
X_2234_ _2236_/A _2234_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_428 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2828__A2 _2910_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_664 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_2165_ _2163_/A _2165_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_656 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_634 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4610__RESET_B _2163_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_325 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3789__B1 _4489_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_509 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_723 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2770__A _4493_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_266 VGND VPWR sky130_fd_sc_hd__decap_8
X_2998_ _2997_/X _3216_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_299 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2764__B2 _4496_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3619_ _3640_/B _3620_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3308__A3 _3307_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_712 VGND VPWR sky130_fd_sc_hd__fill_2
X_4599_ _4220_/Y _3990_/A _2177_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_115_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3106__A _3105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_22 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2945__A _2935_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_111 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4582__D _4582_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4389__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_689 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4244__A2_N _3399_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4351__RESET_B _2473_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_550 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2680__A _2680_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3795__A3 _4491_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_244 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3495__B _3486_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_248 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2755__A1 _2715_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_704 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_428 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3016__A _4357_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2855__A _2855_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_642 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4275__A4 _4213_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4439__RESET_B _2368_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_686 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4492__D _4492_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_656 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_475 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_442 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_667 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3235__A2 _3234_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3970_ _4324_/Q _3960_/B _3970_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_2921_ _2920_/X _2922_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2994__A1 _2908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2590__A _2589_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2852_ _4353_/Q _2851_/X _2852_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_2783_ _2782_/X _2783_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_636 VGND VPWR sky130_fd_sc_hd__fill_2
X_4522_ _3843_/X _4522_/Q _2269_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_4453_ _2631_/X _2804_/A _2351_/X _4450_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_168 VGND VPWR sky130_fd_sc_hd__decap_12
X_3404_ _4240_/B _3386_/X _3412_/A _3405_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_98_520 VGND VPWR sky130_fd_sc_hd__fill_2
X_4384_ _3642_/X _4384_/Q _2434_/X _4551_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2749__B _3820_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_352 VGND VPWR sky130_fd_sc_hd__fill_2
X_3335_ _2895_/X _3335_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3266_ _4330_/Q _3266_/B _3266_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_586 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_547 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_2217_ _2238_/A _2217_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4531__CLK _4539_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2765__A _4495_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_686 VGND VPWR sky130_fd_sc_hd__decap_4
X_3197_ _3045_/X _3196_/X _3114_/X _3209_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_66_483 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_100 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_442 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_667 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_520 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3596__A _3585_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_391 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_586 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2737__A1 _2724_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3934__B1 _2552_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_531 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_402 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_330 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4577__D _4134_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_457 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_428 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4532__RESET_B _2257_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4111__B1 _4026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2675__A _2645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_472 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_450 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_163 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_645 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2825__D _2824_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_70 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2976__A1 _3289_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_391 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_350 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_9 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4404__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3953__B _3417_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_127 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3672__C _3671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4487__D _3787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_683 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_160 VGND VPWR sky130_fd_sc_hd__fill_2
X_3120_ _3071_/A _3120_/B _3023_/Y _3016_/Y _3120_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4554__CLK _4619_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_490 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4102__B1 _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2585__A _2585_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3051_ _3050_/X _3051_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_35_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_689 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_294 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_147 VGND VPWR sky130_fd_sc_hd__decap_6
X_3953_ _4348_/Q _3417_/D _3953_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3884_ _3884_/A _3877_/B _3884_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2967__B2 _2966_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2904_ _2901_/X _2902_/X _2904_/C _2904_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__4483__SET_B _2315_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2835_ _4318_/Q _2831_/X _2834_/X _2835_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4024__B _4024_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3916__B1 _2552_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk_i clkbuf_3_6_0_clk_i/X clkbuf_4_13_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3863__B _3859_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2766_ _4491_/Q _2766_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_8_590 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_606 VGND VPWR sky130_fd_sc_hd__decap_4
X_2697_ _2687_/X _2689_/Y _2694_/X _2696_/X _4447_/D VGND VPWR sky130_fd_sc_hd__a211o_4
X_4505_ _3821_/Y _4505_/Q _2289_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_116 VGND VPWR sky130_fd_sc_hd__decap_4
X_4436_ _4436_/D _2604_/A _2371_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4397__D _3571_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_704 VGND VPWR sky130_fd_sc_hd__fill_2
X_4367_ _3409_/Y _4270_/A _2454_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_661 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_501 VGND VPWR sky130_fd_sc_hd__decap_8
X_3318_ _4376_/Q _2906_/X _2887_/X _3320_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_112_193 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_247 VGND VPWR sky130_fd_sc_hd__fill_2
X_4298_ _3960_/B _4292_/Y _4297_/Y _4618_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3249_ _3243_/X _3251_/A _3247_/X _2917_/B _3248_/X _3249_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XANTENNA__2495__A _2495_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_409 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_114 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2661__C _2659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4215__A _4213_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_350 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4427__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3907__B1 _3906_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_567 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_433 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_422 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_538 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3922__A3 _3920_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_499 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4577__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_309 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3686__A2 _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_523 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_203 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_265 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_287 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_298 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_707 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_100 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_637 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_283 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_434 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2852__B _2851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_136 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2949__A1 _2928_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_158 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_219 VGND VPWR sky130_fd_sc_hd__fill_1
X_2620_ _4510_/Q _2620_/B _2620_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3964__A _3964_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_376 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3913__A3 _3911_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2551_ _3925_/A _2552_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2482_ _2496_/A _2485_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_447 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4454__RESET_B _2350_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4075__A2_N _4565_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4221_ _4595_/Q _2743_/A _4116_/C _2704_/A _2755_/X _4221_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_110_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_320 VGND VPWR sky130_fd_sc_hd__decap_12
X_4152_ _4582_/Q _4153_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3103_ _3102_/X _3103_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4083_ utmi_data_out_o[5] _4082_/X _4083_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_110_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3204__A _3065_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3034_ _3120_/B _3347_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_272 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_412 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4013__A2_N _4012_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_626 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2762__B _2762_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_659 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_467 VGND VPWR sky130_fd_sc_hd__fill_2
X_3936_ _3186_/A _4278_/C _3936_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3867_ _4541_/Q _3859_/B _3867_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3798_ _2601_/X _3785_/X _4494_/Q _4524_/Q _3792_/X _3798_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_2818_ _2818_/A _2799_/A _2818_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3593__B _3593_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2749_ _4501_/Q _3820_/A _3810_/A _4504_/Q _2749_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__3365__A1 _3039_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4201__C _4201_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4419_ _3477_/Y _2900_/A _2392_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_120_439 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_631 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_523 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_239 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3114__A _3011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_22 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4093__A2 _4016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3840__A2 _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_626 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_423 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_99 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3487__C _3486_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4590__D _4590_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_670 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3784__A _3784_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_191 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_417 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_629 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_491 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_504 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_707 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3024__A _3023_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_507 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3959__A _3959_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2863__A _4414_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_389 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_570 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_592 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3678__B _3678_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_423 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2582__B _4552_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_264 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3397__C _3396_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_128 VGND VPWR sky130_fd_sc_hd__decap_4
X_3721_ _2643_/Y _3673_/A _2673_/X _3674_/C _3723_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_9_140 VGND VPWR sky130_fd_sc_hd__decap_8
X_3652_ _3581_/A _3652_/B _3651_/X _3652_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_9_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_184 VGND VPWR sky130_fd_sc_hd__decap_4
X_3583_ _3554_/A _3583_/B _3583_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2603_ _3993_/B _2599_/X _2602_/X _2603_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_115_712 VGND VPWR sky130_fd_sc_hd__decap_12
X_2534_ _2533_/X _2534_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2465_ _2460_/X _2465_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2570__A2 _2554_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2396_ _2396_/A _2399_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_320 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2757__B _2761_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4204_ _2718_/B _2741_/B _2718_/B _4281_/A _4204_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4135_ _2669_/A _4135_/B _4135_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_526 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3869__A _3883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_345 VGND VPWR sky130_fd_sc_hd__decap_3
X_4066_ _4066_/A _4066_/B _4066_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3283__B1 _2928_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2773__A _4492_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_209 VGND VPWR sky130_fd_sc_hd__decap_4
X_3017_ _3015_/X _3016_/Y _4354_/Q _4355_/Q _3017_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_64_581 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_242 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_456 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3919_ _4318_/Q _2585_/A _3919_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_106_701 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4376__RESET_B _2443_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3338__A1 _3334_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4212__B _4211_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2948__A _2948_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_117 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2667__B _2666_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_504 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4615__CLK _4619_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4585__D _4585_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_507 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2683__A _2671_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_570 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3498__B _3498_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3813__A2 _3803_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_423 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_456 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_478 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__C _4105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_489 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_662 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_644 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4122__B _2579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3019__A _3018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_404 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2858__A _3607_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3961__B _4278_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2250_ _2248_/A _2250_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4495__D _4495_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_632 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_172 VGND VPWR sky130_fd_sc_hd__fill_2
X_2181_ _2166_/X _2183_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_77_194 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4057__A2 _4017_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_367 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2593__A _4595_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_581 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3201__B _3198_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_595 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_448 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_314 VGND VPWR sky130_fd_sc_hd__fill_2
X_3704_ _3704_/A _3704_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2953__A2_N _3265_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3635_ outport_data_o[4] _3625_/B _3636_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_108_38 VGND VPWR sky130_fd_sc_hd__fill_2
X_3566_ _3566_/A _3566_/B _3566_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3740__A1 _3671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3740__B2 _3687_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3497_ _3428_/B _3498_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_2517_ _2516_/X _2701_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_2448_ _2449_/A _2448_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_640 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4296__A2 _4292_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2379_ _2379_/A _2379_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_334 VGND VPWR sky130_fd_sc_hd__fill_2
X_4118_ _4115_/X _4116_/X _4117_/X _4118_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_83_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_164 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3599__A _3585_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_4049_ _4566_/Q _4037_/X _4033_/X _4048_/Y _4049_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_71_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3271__A3 _3270_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_215 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_459 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4557__RESET_B _2227_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4220__A2 _4217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_89 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_78 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_380 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_542 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_437 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_120 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3798__A1 _2601_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3302__A _3302_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_592 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3798__B2 _3792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2860__B _2857_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__C _3713_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__C1 _4445_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3972__A _4560_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_60 VGND VPWR sky130_fd_sc_hd__fill_1
X_3420_ _3420_/A _3420_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_3351_ _3359_/A _3347_/Y _3360_/B _3351_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__2588__A _2581_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_234 VGND VPWR sky130_fd_sc_hd__fill_2
X_2302_ _2301_/A _2302_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_680 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_567 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_245 VGND VPWR sky130_fd_sc_hd__decap_6
X_3282_ _3243_/B _2949_/X _3282_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_589 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_481 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_610 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_109 VGND VPWR sky130_fd_sc_hd__fill_2
X_2233_ _2236_/A _2233_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2164_ _2163_/A _2164_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_473 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_101 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3789__A1 _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_581 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4308__A _4247_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3789__B2 _3786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_2997_ _2849_/A _2915_/X _2997_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4043__A _4043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4460__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_339 VGND VPWR sky130_fd_sc_hd__decap_4
X_3618_ _3617_/X _3640_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2498__A _2497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_4598_ _4212_/X _3987_/A _2178_/X _4497_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3549_ _3508_/A _3555_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_103_512 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_223 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_429 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_613 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_507 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_315 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3122__A _3363_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_679 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_540 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2961__A _2922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_370 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2680__B _2679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4391__RESET_B _2426_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_554 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4320__RESET_B _2509_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3776__A1_N _3681_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2755__A2 _2745_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3792__A _3792_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_411 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_38 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_201 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_234 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2201__A _2199_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_23_0_clk_i_A clkbuf_5_22_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_683 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_51 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2855__B _2855_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_473 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_451 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_142 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2970__A1_N _3491_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4333__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3032__A _3015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_679 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4408__RESET_B _2405_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2920_ _4329_/Q _2920_/B _2920_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2871__A _2880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_510 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2994__A2 _2916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4483__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2851_ _2850_/X _2851_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2782_ _2781_/X _2782_/X VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_604 VGND VPWR sky130_fd_sc_hd__fill_2
X_4521_ _3840_/X _4521_/Q _2270_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_125 VGND VPWR sky130_fd_sc_hd__fill_2
X_4452_ _2681_/Y _2785_/C _2352_/X _4450_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_158 VGND VPWR sky130_fd_sc_hd__decap_8
X_3403_ _4267_/A _4240_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_4383_ _3639_/X _2853_/D _2435_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2749__C _3810_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3207__A _3207_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_565 VGND VPWR sky130_fd_sc_hd__fill_1
X_3334_ _3333_/X _3334_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3265_ _3265_/A _3265_/B _3265_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_364 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_504 VGND VPWR sky130_fd_sc_hd__decap_6
X_2216_ _2210_/X _2216_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_54_613 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_676 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_142 VGND VPWR sky130_fd_sc_hd__decap_8
X_3196_ _3031_/X _3360_/A _3196_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_93_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4038__A _4030_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_454 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_156 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3877__A _4545_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2781__A _3707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3596__B _3596_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2737__A2 _2735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3934__A1 _2578_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3934__B2 _3933_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_670 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3117__A _3347_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_554 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2956__A _2917_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_576 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_204 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_248 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4356__CLK _4356_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_99 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4111__B2 _4110_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2675__B _2649_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_440 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4593__D _4593_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_131 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_359 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2691__A _2691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_487 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4501__RESET_B _2293_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_627 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_98 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2976__A2 _2972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_607 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_8 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3672__D _4472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_670 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3689__B1 _2643_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3027__A _4355_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2897__D1 _2872_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2866__A _2866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_513 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_695 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_83 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_72 VGND VPWR sky130_fd_sc_hd__decap_4
X_3050_ _3049_/X _3050_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_82_207 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4102__B2 _4108_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2664__A1 _2691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_638 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_167 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_318 VGND VPWR sky130_fd_sc_hd__fill_1
X_3952_ _4322_/Q _2585_/A _3952_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_16_381 VGND VPWR sky130_fd_sc_hd__fill_2
X_3883_ _3883_/A _3883_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2903_ _3455_/A _3460_/A _3464_/A _3653_/A _2904_/C VGND VPWR sky130_fd_sc_hd__or4_4
X_2834_ inport_data_i[1] inport_accept_o _2834_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3916__B2 _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3916__A1 _2578_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_412 VGND VPWR sky130_fd_sc_hd__fill_2
X_2765_ _4495_/Q _2765_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4504_ _4504_/D _4504_/Q _2290_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2696_ _2696_/A _2696_/B _2695_/X _2696_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_6_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_81 VGND VPWR sky130_fd_sc_hd__fill_2
X_4435_ _4435_/D _2610_/A _2372_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_640 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4379__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4366_ _3405_/Y _4267_/A _2455_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4243__A2_N _3388_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_362 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_513 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2776__A _2771_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3317_ _3317_/A _3316_/Y _3317_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_58_215 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_204 VGND VPWR sky130_fd_sc_hd__fill_2
X_4297_ _2528_/C _3960_/B _2684_/X _4297_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_3248_ _3248_/A _3248_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_462 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_602 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3852__B1 _3851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_473 VGND VPWR sky130_fd_sc_hd__fill_2
X_3179_ _3013_/X _3177_/X _3178_/X _3179_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_27_635 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_432 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_627 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_24 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4215__B _4215_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_362 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2661__D _2660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_671 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_513 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_373 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3907__A1 _3889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_445 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4231__A _2908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4588__D _4181_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_673 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_579 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4096__B1 _4030_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_613 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3843__B1 _3842_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_616 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_446 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3310__A _2986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_649 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2949__A2 _2968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_192 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4020__B1 _4016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4521__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2550_ _2701_/A _2549_/X _2550_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_5_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4141__A _4140_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4498__D _3807_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_572 VGND VPWR sky130_fd_sc_hd__fill_2
X_2481_ _2475_/X _2481_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_459 VGND VPWR sky130_fd_sc_hd__fill_2
X_4220_ _2704_/A _4217_/X _4219_/X _3990_/Y _4207_/X _4220_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_5_594 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3980__A utmi_txready_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_513 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_332 VGND VPWR sky130_fd_sc_hd__decap_12
X_4151_ _4143_/X _4151_/B _4150_/Y _4151_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__2596__A _2596_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_354 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4494__RESET_B _2302_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_3102_ _3007_/X _3038_/Y _4358_/Q _4359_/Q _3102_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4087__B1 _3957_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4082_ _4018_/Y _4081_/X _4018_/Y _4081_/X _4082_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4423__RESET_B _2387_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_270 VGND VPWR sky130_fd_sc_hd__fill_1
X_3033_ _4357_/Q _3360_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3204__B _3122_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2762__C _2762_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3220__A _3108_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_638 VGND VPWR sky130_fd_sc_hd__decap_3
X_3935_ _4320_/Q _2585_/A _3935_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_31_170 VGND VPWR sky130_fd_sc_hd__decap_4
X_3866_ _4532_/Q _3855_/X _3865_/X _3866_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_31_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_3797_ _2601_/X _3785_/X _4493_/Q _2645_/X _3792_/X _3797_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_2817_ _2818_/A _2821_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3593__C _3592_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2748_ _4499_/Q _4498_/Q _2750_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3365__A2 _3364_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_297 VGND VPWR sky130_fd_sc_hd__fill_2
X_4418_ _3474_/Y _4418_/Q _2393_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2679_ _2657_/X _2658_/Y _2678_/X _2679_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_120_407 VGND VPWR sky130_fd_sc_hd__decap_4
X_4349_ _3226_/Y _4349_/Q _2476_/X _4325_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_101_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_410 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3114__B _3369_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4562__SET_B _2221_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_571 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_593 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_435 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_11 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4544__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_231 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_220 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3761__C1 _3760_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4305__A1 _4467_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_520 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_597 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3305__A _3317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4069__B1 _3933_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_376 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_410 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2863__B _2863_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_95 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3678__C _3677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3040__A _4361_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4136__A _4135_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_608 VGND VPWR sky130_fd_sc_hd__fill_2
X_3720_ _3720_/A _3724_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4241__B1 _4266_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_529 VGND VPWR sky130_fd_sc_hd__fill_2
X_3651_ _3522_/A _3646_/Y _3651_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3582_ _3582_/A _3582_/B _3582_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_61_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_2602_ _2601_/X _2602_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_724 VGND VPWR sky130_fd_sc_hd__fill_1
X_2533_ _2532_/X _2533_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_107 VGND VPWR sky130_fd_sc_hd__decap_8
X_2464_ _2460_/X _2464_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2395_ _2391_/A _2395_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4604__RESET_B _2171_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4203_ _2516_/X _4202_/Y _4143_/X _4593_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_3_82 VGND VPWR sky130_fd_sc_hd__fill_2
X_4134_ _2736_/X _4132_/X _4134_/C _4134_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3215__A _4349_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_473 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4417__CLK _4410_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3807__B1 _3806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_549 VGND VPWR sky130_fd_sc_hd__fill_2
X_4065_ _4066_/A _4066_/B _4065_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3283__B2 _3277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3283__A1 _3280_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3016_ _4357_/Q _3016_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_64_593 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_221 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4567__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4046__A _4046_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_287 VGND VPWR sky130_fd_sc_hd__decap_8
X_3918_ _4562_/Q _3918_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3849_ _4533_/Q _3844_/X _3849_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2794__B1 _2639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_7 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3338__A2 _3337_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3743__C1 _3742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_306 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4212__C _4212_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_716 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_267 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_215 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_321 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4345__RESET_B _2480_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_248 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_451 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_207 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2964__A _2955_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2683__B _2631_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_251 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3498__C _3498_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_593 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_76 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_276 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4223__B1 _4602_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_49 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_634 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_144 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_122 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2204__A _2206_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_73 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2858__B _2858_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_140 VGND VPWR sky130_fd_sc_hd__decap_4
X_2180_ _2177_/A _2180_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3035__A _3359_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_685 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_151 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4027__A2_N _4026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_184 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2874__A _2874_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3201__C _3200_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4214__B1 _4213_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_287 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_416 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_326 VGND VPWR sky130_fd_sc_hd__fill_1
X_3703_ _3702_/A _3701_/X _3720_/A _3702_/Y _3705_/B VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_119_359 VGND VPWR sky130_fd_sc_hd__decap_3
X_3634_ _3634_/A _3620_/B _3634_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3725__C1 _3724_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_17 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_3565_ _3555_/A _3565_/B _3564_/X _3565_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_115_576 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3740__A2 _3687_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3496_ _3504_/A _3494_/Y _3495_/X _4425_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_88_416 VGND VPWR sky130_fd_sc_hd__decap_12
X_2516_ _2696_/A _2516_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_2447_ _2449_/A _2447_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_259 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_248 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_237 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_652 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2700__B1 _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2378_ _2379_/A _2378_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_696 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_313 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2784__A _2784_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4117_ _3987_/Y _4602_/Q _3987_/A _3999_/Y _4117_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3599__B _3597_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4048_ _4048_/A _4073_/A _4048_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_17_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_582 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_216 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_541 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_703 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_238 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_714 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2767__B1 _4608_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4220__A3 _4219_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4597__RESET_B _2179_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_471 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3716__C1 _3715_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_532 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4526__RESET_B _2264_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_648 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4596__D _4208_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_43 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_281 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_493 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2694__A _2694_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_633 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_335 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_305 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_64 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3302__B _3246_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3798__A2 _3785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_287 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2860__C _2860_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_393 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_235 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__B1 _2628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3675__D _3711_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_392 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2869__A _4379_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_703 VGND VPWR sky130_fd_sc_hd__fill_2
X_3350_ _3347_/A _3347_/B _3350_/C _3325_/X _3360_/B VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__2588__B _2587_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3183__B1 _3240_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2301_ _2301_/A _2301_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3281_ _2928_/A _3275_/B _3281_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_279 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_302 VGND VPWR sky130_fd_sc_hd__fill_1
X_2232_ _2236_/A _2232_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_24_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2163_ _2163_/A _2163_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_463 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_560 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_508 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_113 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_316 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4308__B _2707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_669 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3789__A2 _3782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_393 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_112 VGND VPWR sky130_fd_sc_hd__fill_2
X_2996_ _2996_/A _2908_/X _2995_/Y _2996_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_119_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4605__CLK _4619_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4043__B _4039_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_156 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_189 VGND VPWR sky130_fd_sc_hd__fill_2
X_3617_ _3616_/X _3617_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2779__A _2778_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4597_ _4209_/X _3984_/A _2179_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3548_ _3545_/A _3546_/Y _3547_/X _4407_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_103_535 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_502 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106 VGND VPWR sky130_fd_sc_hd__decap_12
X_3479_ _3510_/A _3479_/B _3480_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_103_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_460 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_121 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3403__A _4267_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_688 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_379 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_496 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_625 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2809__B1_N _2808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2988__B1 _3460_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_585 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_40 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4234__A _4234_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_55 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2689__A _3713_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4360__RESET_B _2462_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_423 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_343 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4114__C1 _4113_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_290 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_695 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2855__C _3582_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_74 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3313__A _3317_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_27_0_clk_i_A clkbuf_4_13_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_625 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_146 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2871__B _2871_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_585 VGND VPWR sky130_fd_sc_hd__fill_1
X_2850_ _2905_/A _2850_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_43_382 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4144__A _4144_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_596 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2967__A2_N _2966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _3707_/A _2633_/X _2781_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4448__RESET_B _2357_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3983__A _2701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4520_ _3838_/X _4520_/Q _2271_/X _4519_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_649 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_137 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_115 VGND VPWR sky130_fd_sc_hd__fill_2
X_4451_ _2671_/D _2784_/A _2354_/X _4509_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2599__A _3994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_148 VGND VPWR sky130_fd_sc_hd__fill_1
X_3402_ _2858_/B _3398_/B _3402_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3156__B1 _3066_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4382_ _3636_/X _3634_/A _2436_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2749__D _4504_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3207__B _3199_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3333_ _3330_/X _3332_/X _3333_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3264_ _3268_/A _3264_/B _4329_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_39_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_387 VGND VPWR sky130_fd_sc_hd__decap_8
X_2215_ _2210_/X _2215_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_655 VGND VPWR sky130_fd_sc_hd__fill_2
X_3195_ _3366_/A _2916_/Y _4347_/Q _3195_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_38_154 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3223__A _3085_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_411 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_466 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_349 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3877__B _3877_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2781__B _2633_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3596__C _3595_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_680 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4054__A _4073_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_511 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3893__A utmi_data_in_i[0] VGND VPWR sky130_fd_sc_hd__diode_2
X_2979_ _2979_/A _2979_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_22_599 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_209 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3934__A2 _3932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2302__A _2301_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3147__B1 _3146_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_118 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3117__B _3035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_376 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2956__B _2917_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_290 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4229__A _4278_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3133__A _2996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_636 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3682__A2_N _3675_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2972__A _2972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_146 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2691__B _2691_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_499 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_691 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3697__A2_N _3696_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4541__RESET_B _2246_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3689__A1 _4520_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3689__B2 _2641_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_264 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2212__A _2210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_181 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2897__C1 _2876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_80 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_503 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_184 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2866__B _2863_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_536 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_709 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4139__A _4138_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3043__A _3031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4450__CLK _4450_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2664__A2 _2670_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_444 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_658 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3978__A _3978_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_628 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_105 VGND VPWR sky130_fd_sc_hd__decap_8
X_3951_ _3950_/X utmi_data_out_o[4] VGND VPWR sky130_fd_sc_hd__buf_1
X_2902_ _3488_/A _3491_/A _3494_/A _2902_/D _2902_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_50_116 VGND VPWR sky130_fd_sc_hd__decap_8
X_3882_ _4539_/Q _3869_/X _3881_/X _3882_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_91_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_330 VGND VPWR sky130_fd_sc_hd__fill_2
X_2833_ _4317_/Q _2831_/X _2832_/X _2833_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_2764_ _4234_/A _4496_/Q _4234_/A _4496_/Q _2764_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__3377__B1 _3376_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3916__A2 _3914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4503_ _3817_/Y _4503_/Q _2291_/X _4450_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_581 VGND VPWR sky130_fd_sc_hd__fill_2
X_2695_ _2694_/A _3717_/A _2804_/A _2695_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3130__A1_N _3029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_4434_ _2617_/X _4050_/A _2373_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
X_4365_ _3401_/Y _3399_/A _2456_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_685 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_3316_ _3251_/A _3314_/X _3315_/X _3314_/A _3248_/A _3316_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_100_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2776__B _2772_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4296_ _2725_/Y _4292_/Y _4295_/Y _4296_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3247_ _2917_/B _3266_/B _3247_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_86_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_379 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3852__A1 _2659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_260 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_485 VGND VPWR sky130_fd_sc_hd__decap_3
X_3178_ _3058_/X _3047_/X _3178_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_66_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_647 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_488 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_14 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_308 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_319 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_499 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_691 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_7_0_clk_i clkbuf_4_7_0_clk_i/A clkbuf_4_7_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_50_683 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_503 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3907__A2 _3897_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3368__B1 _3367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4231__B _3238_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3128__A _3123_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4323__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3728__A1_N _3674_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_514 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4473__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_396 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2984__A1_N _3451_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_249 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4096__A1 _4093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3843__A1 _3685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_580 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3310__B _3246_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_661 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2207__A _2206_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4020__B2 _4019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3038__A _4360_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_562 VGND VPWR sky130_fd_sc_hd__decap_8
X_2480_ _2475_/X _2480_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_90 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2877__A _2876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3980__B _3980_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4150_ _4153_/A _4147_/C _4150_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_68_536 VGND VPWR sky130_fd_sc_hd__fill_2
X_3101_ _3221_/A _3171_/A _3190_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_95_344 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4087__B2 _4007_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4081_ _3949_/Y _4566_/Q _3949_/Y _4566_/Q _4081_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_539 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_528 VGND VPWR sky130_fd_sc_hd__fill_2
X_3032_ _3015_/X _3359_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3501__A _4410_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_550 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4463__RESET_B _2340_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2762__D _2761_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3220__B _3137_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3934_ _2578_/X _3932_/X _2552_/A _3933_/Y utmi_data_out_o[2] VGND VPWR sky130_fd_sc_hd__o22a_4
X_3865_ _4540_/Q _3859_/B _3865_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_32_672 VGND VPWR sky130_fd_sc_hd__fill_2
X_2816_ _2815_/X _2825_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4346__CLK _4342_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3796_ _2684_/X _3785_/X _4492_/Q _3685_/X _3792_/X _4492_/D VGND VPWR sky130_fd_sc_hd__a32o_4
X_2747_ _4502_/Q _3814_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_254 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_416 VGND VPWR sky130_fd_sc_hd__decap_8
X_2678_ _2673_/X _2674_/Y _2661_/X _2654_/B _2677_/Y _2678_/X VGND VPWR sky130_fd_sc_hd__o32a_4
X_4417_ _3526_/Y _2863_/B _2394_/X _4410_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4496__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2787__A _2786_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_600 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_503 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_110 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_536 VGND VPWR sky130_fd_sc_hd__decap_8
X_4348_ _3213_/X _4348_/Q _2477_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_100_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_569 VGND VPWR sky130_fd_sc_hd__fill_2
X_4279_ _4277_/Y _4278_/X _4280_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_101_699 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_400 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3114__C _3046_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_293 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_13 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_422 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_433 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3411__A _4392_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_466 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_469 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_672 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_491 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_344 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4242__A _4242_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_315 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_366 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_359 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4599__D _4220_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3761__B1 _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4305__A2 _2782_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_333 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3305__B _3304_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_325 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_399 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_388 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4069__B2 _4022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_369 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_701 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_414 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4369__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3040__B _3038_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_469 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_447 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4241__B2 _4267_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_288 VGND VPWR sky130_fd_sc_hd__decap_4
X_3650_ _4376_/Q _3646_/Y _3652_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4152__A _4582_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_153 VGND VPWR sky130_fd_sc_hd__fill_2
X_3581_ _3581_/A _3579_/Y _3581_/C _3581_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_2601_ _2601_/A _2601_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3752__B1 _3683_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2532_ _4489_/Q _4488_/Q _2531_/Y _2532_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_54_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_246 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_2463_ _2460_/X _2463_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4202_ _4185_/Y _4194_/Y _4198_/Y _4202_/D _4202_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__2400__A _2399_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2394_ _2391_/A _2394_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_4133_ _2575_/A _4127_/X _3979_/X _4134_/C VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_29_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_675 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_377 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_366 VGND VPWR sky130_fd_sc_hd__fill_2
X_4064_ _4562_/Q _4563_/Q _3918_/Y _3933_/Y _4066_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_28_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_496 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_196 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_336 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3807__A1 _2643_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3015_ _4356_/Q _3015_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3283__A2 _3281_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_561 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4046__B _4073_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_414 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2794__A1 _2635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_3917_ _3916_/X utmi_data_out_o[0] VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_491 VGND VPWR sky130_fd_sc_hd__decap_4
X_3848_ _4524_/Q _3841_/X _3847_/X _3848_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3991__B1 _3937_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4062__A _4073_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_26 VGND VPWR sky130_fd_sc_hd__fill_1
X_3779_ _3724_/A _3674_/D _2687_/X _3778_/X _3779_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_118_552 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3743__B1 _3719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_596 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3406__A _3607_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2310__A _2324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2964__B _2957_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_196 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4385__RESET_B _2433_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_78 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_56 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4511__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_358 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2683__C _2682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_550 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4237__A _4612_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3141__A _3138_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_62 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_263 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_55 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4223__A1 _2704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4223__B2 _2706_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_4_0_clk_i clkbuf_2_2_0_clk_i/X clkbuf_4_9_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_141 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3982__B1 _3912_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_541 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_112 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3734__B1 _3702_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_167 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_41 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2858__C _4393_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_384 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2220__A _2217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_642 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3035__B _3360_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_561 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3051__A _3050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4147__A _4143_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_520 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_712 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_285 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3986__A _2701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_575 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4214__A1 _2534_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_3702_ _3702_/A _3701_/X _3702_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3973__B1 _2581_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3633_ _3662_/A _3633_/B _3632_/X _3633_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3725__B1 _3719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_3564_ _3506_/A _3582_/B _3564_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_544 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_717 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_706 VGND VPWR sky130_fd_sc_hd__decap_4
X_3495_ _3554_/A _3486_/B _3495_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_2515_ _2628_/C _2696_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_2446_ _2425_/A _2449_/A VGND VPWR sky130_fd_sc_hd__buf_1
Xclkbuf_5_6_0_clk_i clkbuf_4_3_0_clk_i/X _4619_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3226__A _3397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_260 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4534__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_612 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2700__B2 _2699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2700__A1 _4510_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2377_ _2379_/A _2377_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4116_ _4116_/A _3984_/Y _4116_/C _4116_/D _4116_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_83_111 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2784__B _4449_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3599__C _3598_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2768__A1_N _4242_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VPWR sky130_fd_sc_hd__fill_2
X_4047_ _4565_/Q _4037_/X _4033_/X _4046_/Y _4565_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_83_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_206 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_553 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_244 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_439 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2305__A _2306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2767__B2 _2766_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_450 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_483 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3716__B1 _3704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_605 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_627 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_555 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_409 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2975__A _2933_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2694__B _2694_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_196 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_347 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_72 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_200 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3798__A3 _4494_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_203 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_704 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_715 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_64 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_597 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_299 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2215__A _2210_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2758__A1 _4050_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4407__CLK _4407_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_432 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_461 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_308 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_476 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_498 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3183__A1 _3928_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_225 VGND VPWR sky130_fd_sc_hd__fill_2
X_2300_ _2301_/A _2300_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3280_ _3251_/A _3280_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3046__A _3007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4557__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2231_ _2238_/A _2236_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_78_450 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2885__A _4376_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2162_ _2163_/A _2162_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_17_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_615 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_656 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_369 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_648 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4308__C _4307_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3789__A3 _3790_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_564 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_715 VGND VPWR sky130_fd_sc_hd__decap_8
X_2995_ _2916_/Y _2993_/X _2994_/X _2995_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_9_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3946__B1 _2604_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_82 VGND VPWR sky130_fd_sc_hd__fill_2
X_3616_ _3426_/Y _3427_/B _3528_/C _3498_/C _3616_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_5_1_0_clk_i_A clkbuf_5_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4596_ _4208_/X _3978_/A _2180_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3547_ _3547_/A _3544_/B _3547_/X VGND VPWR sky130_fd_sc_hd__and2_4
Xclkbuf_5_29_0_clk_i clkbuf_5_29_0_clk_i/A _4423_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_1_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_619 VGND VPWR sky130_fd_sc_hd__decap_4
X_3478_ _4420_/Q _3478_/B _3478_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4123__B1 _2608_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2429_ _2431_/A _2429_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_314 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_133 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_24 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2988__B2 _2987_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_383 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_247 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_67 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4026__A2_N _4025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2689__B _2689_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4250__A _4249_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_446 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4400__D _3581_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4114__B1 _4033_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_355 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_601 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_641 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_591 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2855__D _4400_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3313__B _3312_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4472__SET_B _2328_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_103 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_564 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_681 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_394 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_523 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ _2696_/B _2779_/Y _2780_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3983__B _3983_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_clk_i clkbuf_2_1_0_clk_i/A clkbuf_3_3_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_291 VGND VPWR sky130_fd_sc_hd__fill_2
X_4450_ _4450_/D _4450_/Q _2355_/X _4450_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4488__RESET_B _2309_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_262 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4160__A _4160_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2599__B _4437_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4417__RESET_B _2394_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4381_ _3633_/X _3331_/D _2437_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3401_ _3398_/Y _3400_/X _3401_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3156__B2 _3036_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_30_0_clk_i clkbuf_5_30_0_clk_i/A _4410_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_3332_ _4378_/Q _2869_/Y _3332_/C _2872_/B _3332_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_112_322 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_545 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_707 VGND VPWR sky130_fd_sc_hd__decap_12
X_3263_ _3251_/X _3261_/X _3262_/X _4329_/Q _3248_/X _3264_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_112_377 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3504__A _3504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_239 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_280 VGND VPWR sky130_fd_sc_hd__decap_3
X_3194_ _2850_/X _3366_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_2214_ _2210_/X _2214_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3223__B _3223_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_648 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_478 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_383 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_16 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4054__B _4054_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3893__B _3895_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2978_ _2950_/Y _2971_/X _2974_/Y _2978_/D _2978_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_107_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_138 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3147__A1 _3041_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_59 VGND VPWR sky130_fd_sc_hd__decap_3
X_4579_ _4142_/X _4135_/B _2200_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_438 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3117__C _3014_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_589 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_707 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clk_i clkbuf_4_3_0_clk_i/A clkbuf_4_3_0_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3414__A _3414_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4229__B _4278_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3133__B _3133_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4245__A _4240_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_342 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_364 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4032__C1 _4031_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4581__RESET_B _2198_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_672 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3689__A2 _2657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4510__RESET_B _2283_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_193 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2897__B1 _3331_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_664 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2866__C _2864_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_228 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3324__A _2913_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3043__B _3105_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_489 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4155__A _4143_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3950_ _2578_/X _3948_/X _2552_/A _3949_/Y _3950_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3074__B1 _3065_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2901_ _4427_/Q _4428_/Q _4429_/Q _3451_/A _2901_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_3881_ _4547_/Q _3877_/B _3881_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3994__A _3994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2832_ inport_data_i[0] inport_accept_o _2832_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_31_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_2763_ _2763_/A _2763_/B _2763_/C _2725_/Y outport_valid_o VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__3377__A1 _3375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2403__A _2396_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_4502_ _3815_/Y _4502_/Q _2292_/X _4450_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_469 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_458 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_447 VGND VPWR sky130_fd_sc_hd__decap_4
X_2694_ _2694_/A _2694_/B _2694_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4433_ _3467_/Y _3464_/A _2375_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4364_ _4364_/D _4260_/A _2457_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_653 VGND VPWR sky130_fd_sc_hd__fill_2
X_3315_ _3253_/A _2991_/B _3315_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4295_ _2524_/C _2725_/Y _4247_/A _4295_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__2776__C _2776_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3246_ _3246_/A _3266_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3234__A _2913_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_196 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3127__A2_N _3103_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3757__A2_N _3668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_581 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3852__A2 _3841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_412 VGND VPWR sky130_fd_sc_hd__decap_4
X_3177_ _3110_/C _3363_/A _3097_/X _3177_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_27_615 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_456 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4065__A _4066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_106 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4058__A1_N _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_48 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_14 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4339__RESET_B _2487_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3368__A1 _2851_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_47 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2313__A _2314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3409__A _3406_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4231__C _4231_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3128__B _3124_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_642 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_331 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4618__CLK _4619_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_257 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_11 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3144__A _4358_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_22 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4096__A2 _4095_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_272 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3843__A2 _3841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_592 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_445 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_478 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_94 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3056__B1 _3055_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_695 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_70 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_183 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3319__A _3319_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2223__A _2217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_439 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_504 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_548 VGND VPWR sky130_fd_sc_hd__decap_4
X_3100_ _3227_/D _3084_/A _3171_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3054__A _3381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3989__A _2701_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4080_ _3931_/A _4056_/X _4050_/X _4079_/Y _4571_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_95_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_518 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2893__A _2880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3295__B1 _3293_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_209 VGND VPWR sky130_fd_sc_hd__fill_2
X_3031_ _4354_/Q _3031_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_76_592 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_445 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3501__B _3512_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_540 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_595 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_584 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_437 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_681 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3220__C _3220_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3933_ _4563_/Q _3933_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_640 VGND VPWR sky130_fd_sc_hd__fill_1
X_3864_ _4531_/Q _3855_/X _3863_/X _3864_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4432__RESET_B _2376_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2815_ _2788_/A _2809_/X _2811_/X _2814_/Y _2815_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_118_723 VGND VPWR sky130_fd_sc_hd__fill_2
X_3795_ _2684_/X _3782_/X _4491_/Q _2657_/X _3792_/X _4491_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__3229__A _4350_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_211 VGND VPWR sky130_fd_sc_hd__decap_8
X_2746_ _4219_/A _4469_/Q _4282_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_2677_ _2676_/X _2677_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3681__A2_N _4474_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4416_ _3523_/Y _2866_/A _2395_/X _4410_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_105_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_472 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_150 VGND VPWR sky130_fd_sc_hd__decap_3
X_4347_ _3203_/Y _4347_/Q _2478_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_494 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_634 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_345 VGND VPWR sky130_fd_sc_hd__fill_1
X_4278_ _2537_/X _2730_/D _4278_/C _4278_/D _4278_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_86_389 VGND VPWR sky130_fd_sc_hd__decap_4
X_3229_ _4350_/Q _3229_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3114__D _3375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3411__B _3398_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_618 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2308__A _2306_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_640 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_684 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_200 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3139__A _3059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3761__A1 _3726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2978__A _2950_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4440__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_544 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_472 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_345 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4590__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_367 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_0_0_clk_i clkbuf_2_0_0_clk_i/X clkbuf_4_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_92_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_31 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3602__A _3585_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_434 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_562 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_584 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_713 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2218__A _2217_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3040__C _3039_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_481 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_110 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3049__A _3350_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_3580_ _3522_/A _3583_/B _3581_/C VGND VPWR sky130_fd_sc_hd__and2_4
X_2600_ _2628_/C _2601_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_42_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3752__B2 _3690_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3752__A1 _3683_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2531_ _2524_/X _2531_/B _2528_/X _2531_/D _2531_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__2888__A _3392_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_258 VGND VPWR sky130_fd_sc_hd__decap_12
X_2462_ _2460_/X _2462_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_47_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_393 VGND VPWR sky130_fd_sc_hd__fill_2
X_4201_ _4201_/A _4199_/X _4201_/C _4592_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_2393_ _2391_/A _2393_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_122_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_62 VGND VPWR sky130_fd_sc_hd__decap_3
X_4132_ _3993_/B _4131_/X _4132_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_110_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_153 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_710 VGND VPWR sky130_fd_sc_hd__decap_12
X_4063_ _4568_/Q _4056_/X _4050_/X _4062_/Y _4063_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_3_95 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3512__A _4413_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3807__A2 _3803_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3014_ _3013_/X _3014_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_83_359 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3283__A3 _3282_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_426 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_234 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4613__RESET_B _2160_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_459 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_2_0_clk_i clkbuf_5_3_0_clk_i/A _4446_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_3916_ _2578_/X _3914_/Y _2552_/A _3915_/Y _3916_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3847_ _4532_/Q _3844_/X _3847_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4463__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2794__A2 _2790_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3991__B2 _3981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3991__A1 _3990_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4062__B _4062_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_654 VGND VPWR sky130_fd_sc_hd__decap_4
X_3778_ _3698_/Y _3776_/X _3777_/Y _3778_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_118_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_575 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3743__A1 _3726_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2729_ _3812_/A _4505_/Q _2729_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_105_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_621 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3406__B _3398_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_35 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3259__B1 _4328_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2964__C _2960_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3422__A _4372_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_348 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_337 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2683__D _2681_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3141__B _3188_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_381 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_532 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4354__RESET_B _2470_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_459 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__A _4253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_267 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4223__A2 _2733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_407 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_632 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_603 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_654 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3982__B2 _3981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3982__A1 _4116_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4403__D _4403_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_520 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3734__B2 _3680_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3734__A1 _3679_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_575 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_407 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2501__A _2497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_418 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2858__D _4392_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3035__C _3347_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_635 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3332__A _4378_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4336__CLK _4334_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_7 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_679 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4147__B _4147_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_90 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_264 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4486__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_543 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_297 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3986__B _3986_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_587 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4214__A2 _2714_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4163__A _4143_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3701_ _3681_/X _3700_/X _3681_/X _3700_/X _3701_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3973__A1 _2605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3973__B2 _3972_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3632_ outport_data_o[3] _3625_/B _3632_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3725__A1 _3708_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_clk_i_A clkbuf_4_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3507__A _3504_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3563_ _3563_/A _3566_/B _3565_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_567 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2411__A _2411_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3494_ _3494_/A _3479_/B _3494_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_88_407 VGND VPWR sky130_fd_sc_hd__decap_6
X_2514_ _4620_/D _2628_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_2445_ _2443_/A _2445_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3226__B _3216_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2376_ _2379_/A _2376_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2700__A2 _2810_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_687 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_665 VGND VPWR sky130_fd_sc_hd__fill_2
X_4115_ _3990_/Y _4603_/Q _3990_/A _4002_/Y _4115_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_110_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3242__A _3265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_186 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2784__C _2696_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_294 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VPWR sky130_fd_sc_hd__decap_3
X_4046_ _4046_/A _4073_/A _4046_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_25_724 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_25_0_clk_i clkbuf_5_25_0_clk_i/A _4551_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_212 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_229 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_256 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4073__A _4073_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3716__A1 _3708_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_512 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3417__A _2763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_567 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2321__A _2318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_418 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_12 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_559 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4241__A2_N _3388_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4359__CLK _4334_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_112 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4248__A _2696_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4535__RESET_B _2254_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_359 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_189 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2991__A _3464_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_381 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_595 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_384 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3404__B1 _3412_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__A2 _4443_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_259 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_473 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_444 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3327__A _3559_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2231__A _2238_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3183__A2 _2999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_215 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_661 VGND VPWR sky130_fd_sc_hd__fill_2
X_2230_ _2228_/A _2230_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_410 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_123 VGND VPWR sky130_fd_sc_hd__decap_8
X_2161_ _2163_/A _2161_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_326 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4158__A _4187_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3062__A _3061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_668 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_348 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_476 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_329 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3997__A _3994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_690 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2406__A _2408_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2994_ _2908_/C _2916_/Y _2850_/X _2994_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_21_226 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3946__A1 _2581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3946__B2 _4557_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_29 VGND VPWR sky130_fd_sc_hd__decap_4
X_3615_ _3612_/A _3613_/X _3615_/C _4393_/D VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3237__A _4342_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4595_ _4212_/C _4595_/Q _2182_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3546_ _4407_/Q _3543_/B _3546_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4501__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_716 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_3477_ _3483_/A _3475_/Y _3477_/C _3477_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4123__A1 _2577_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_5_0_clk_i_A clkbuf_5_4_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2428_ _2431_/A _2428_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_602 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3882__B1 _3881_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_646 VGND VPWR sky130_fd_sc_hd__decap_4
X_2359_ _2358_/A _2359_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_465 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_318 VGND VPWR sky130_fd_sc_hd__fill_2
X_4029_ _3994_/A _2581_/X _4029_/C _4029_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_71_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_521 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2316__A _2314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_97 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3231__B1_N _3230_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4250__B _4250_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_51 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4568__SET_B _2214_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2986__A _2986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4114__A1 _3974_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_664 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_443 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_432 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_134 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_329 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3610__A _4392_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_137 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_373 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2226__A _2228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_91 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_7 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4524__CLK _4539_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_241 VGND VPWR sky130_fd_sc_hd__decap_3
X_4380_ _3629_/X _2880_/A _2438_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2767__A1_N _4612_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3400_ _3399_/Y _3398_/B _3412_/A _3400_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_3331_ _4376_/Q _4375_/Q _2893_/Y _3331_/D _3332_/C VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_98_557 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2896__A _2896_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3262_ _4329_/Q _3266_/B _3262_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_568 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_719 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4457__RESET_B _2347_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3504__B _3504_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_635 VGND VPWR sky130_fd_sc_hd__decap_4
X_2213_ _2210_/X _2213_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3193_ _2996_/A _3186_/X _3193_/C _3193_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3864__B1 _3863_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_432 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_487 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_605 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_318 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_19 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3520__A _3514_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4054__C _4053_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_568 VGND VPWR sky130_fd_sc_hd__fill_2
X_2977_ _4427_/Q _2976_/X _4427_/Q _2976_/X _2978_/D VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_116_640 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4501__D _3813_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3147__A2 _3151_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_502 VGND VPWR sky130_fd_sc_hd__fill_1
X_4578_ _4129_/Y _2606_/C _2201_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3529_ _3544_/B _3543_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_101 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4229__C _2730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_134 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3133__C _3133_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_616 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_318 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3430__A _3430_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_690 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4245__B _4241_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_310 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4226__A1_N _4207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4547__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_557 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4032__B1 _4030_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4261__A _4265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_712 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_701 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4411__D _3507_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_640 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_244 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_695 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_684 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3605__A _3585_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2897__A1 _4379_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_288 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_676 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_131 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4550__RESET_B _2235_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2866__D _2865_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3324__B _3322_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3846__B1 _3845_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_421 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3043__C _3015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_700 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_413 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_476 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3340__A _3559_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_159 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4155__B _4153_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2900_ _2900_/A _4420_/Q _4421_/Q _2900_/D _2900_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_90_276 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3074__B2 _3073_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_310 VGND VPWR sky130_fd_sc_hd__fill_2
X_3880_ _4538_/Q _3869_/X _3879_/X _4538_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_43_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3994__B _3994_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2831_ _2829_/A _2831_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4023__B1 _3969_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3377__A2 _3369_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2762_ _2757_/X _2762_/B _2762_/C _2761_/X _2762_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4171__A _4197_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4501_ _3813_/Y _4501_/Q _2293_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_2693_ _3720_/A _2691_/X _2692_/Y _2694_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
X_4432_ _3463_/Y _3460_/A _2376_/X _4418_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4321__D _2841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4087__A2_N _4007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3515__A _4414_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_321 VGND VPWR sky130_fd_sc_hd__decap_12
X_4363_ _3393_/Y _4257_/A _2458_/X _4380_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_112_131 VGND VPWR sky130_fd_sc_hd__fill_2
X_3314_ _3314_/A _3246_/A _3314_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4294_ _3657_/D _4292_/Y _4293_/Y _4616_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__4010__A2_N _4009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2776__D _2775_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3245_ _3241_/A _3246_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_39_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_571 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_3176_ _3176_/A _3073_/Y _3176_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_27_627 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3250__A _3268_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_424 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_619 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_16 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4065__B _4066_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_16 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_118 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_13_0_clk_i_A clkbuf_4_6_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4014__B1 utmi_data_out_o[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_354 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_365 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3368__A2 _3365_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_538 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3409__B _3409_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_459 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4231__D _2911_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4379__RESET_B _2440_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3128__C _3125_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_715 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_492 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3425__A _3528_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_538 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_527 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3144__B _3010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3828__B1 _4514_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4256__A _4232_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_413 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3160__A _3137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3056__A1 _3085_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4406__D _3545_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_682 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_162 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_82 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2504__A _2504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_358 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3319__B _3320_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4103__A1_N _4100_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_542 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3335__A _2895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_602 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3054__B _3038_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3819__B1 _3818_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3295__A1 _3280_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3295__B2 _3277_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_262 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3989__B _3988_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3030_ _3029_/X _3085_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_63_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4166__A _4164_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_619 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3070__A _3069_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4244__B1 _4610_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4316__D _2848_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3220__D _3219_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_170 VGND VPWR sky130_fd_sc_hd__decap_12
X_3932_ _2571_/X _3930_/Y _2610_/Y _4041_/A _3932_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3863_ _4539_/Q _3859_/B _3863_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2414__A _2411_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2814_ _2803_/A _2812_/Y _2813_/X _2814_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_32_696 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3755__C1 _3754_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3794_ _2684_/X _3782_/X _4490_/Q _2673_/X _3792_/X _3794_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_117_223 VGND VPWR sky130_fd_sc_hd__fill_2
X_2745_ _4219_/A _2548_/Y _4469_/Q _2745_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_117_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_2676_ _2675_/X _2676_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4415_ _4415_/D _2864_/D _2397_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4401__RESET_B _2413_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_663 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_652 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3245__A _3241_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4346_ _3193_/Y _4346_/Q _2479_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_86_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_657 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4392__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_4277_ _4615_/Q _4277_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3228_ _3228_/A _3227_/X _3228_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_36_26 VGND VPWR sky130_fd_sc_hd__fill_1
X_3159_ _3148_/X _3153_/X _3158_/X _3119_/X _3160_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_82_563 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4235__B1 _4232_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_298 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2797__B1 _4508_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2324__A _2324_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_471 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_713 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2549__B1 _4468_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3139__B _3150_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3761__A2 _3715_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2978__B _2971_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_589 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_578 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3173__A2_N _3172_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3602__B _3602_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_541 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_574 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_265 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4226__B1 _4603_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3040__D _4359_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_663 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2234__A _2236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3049__B _3016_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_1_0_clk_i_A clkbuf_2_0_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3752__A2 _3690_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2530_ _2522_/X _2525_/X _2530_/C _2531_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_114_215 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2960__B1 _4420_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2461_ _2460_/X _2461_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4200_ _4198_/Y _4199_/B _4201_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3065__A _3039_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2392_ _2391_/A _2392_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_324 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_74 VGND VPWR sky130_fd_sc_hd__fill_2
X_4131_ _2562_/X _4130_/X _2587_/Y _4118_/X _4131_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_96_688 VGND VPWR sky130_fd_sc_hd__fill_2
X_4062_ _4073_/A _4062_/B _4061_/X _4062_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3512__B _3512_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_582 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_722 VGND VPWR sky130_fd_sc_hd__decap_3
X_3013_ _3012_/X _3013_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__2409__A _2408_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_254 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4217__B1 _4278_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_393 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2950__A2_N _2949_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_257 VGND VPWR sky130_fd_sc_hd__decap_8
X_3915_ _4561_/Q _3915_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__4608__CLK _4460_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_633 VGND VPWR sky130_fd_sc_hd__fill_2
X_3846_ _2645_/X _3841_/X _3845_/X _3846_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__3991__A2 _3979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4062__C _4061_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3777_ _3698_/Y _3776_/X _3720_/A _3777_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_118_532 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_699 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3743__A2 _3709_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2728_ _4500_/Q _3810_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_105_259 VGND VPWR sky130_fd_sc_hd__fill_2
X_2659_ _4526_/Q _2659_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xclkbuf_5_21_0_clk_i clkbuf_5_21_0_clk_i/A _4356_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_87_611 VGND VPWR sky130_fd_sc_hd__fill_2
X_4329_ _4329_/D _4329_/Q _2499_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_432 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_335 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3259__A1 _3251_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_305 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_700 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3259__B2 _3248_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_498 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_476 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2964__D _2963_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3422__B _3415_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2319__A _2318_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_24 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3141__C _3141_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_405 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4208__B1 _3978_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_287 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4223__A3 _2754_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_460 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_471 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4394__RESET_B _2421_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_666 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3982__A2 _3979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2989__A _3314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4323__RESET_B _2506_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_648 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_677 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3734__A2 _4472_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3195__B1 _4347_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_50 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_587 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_54 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_320 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_292 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3613__A _4393_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_677 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_176 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3332__B _2869_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_349 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2229__A _2228_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4147__C _4147_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_243 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_500 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_276 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_235 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_408 VGND VPWR sky130_fd_sc_hd__fill_2
X_3700_ _3682_/X _3699_/X _3682_/X _3699_/X _3700_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4163__B _4161_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_318 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3973__A2 _3970_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3631_ _3331_/D _3620_/B _3633_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3725__A2 _3668_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3562_ _3555_/A _3562_/B _3561_/X _3562_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3507__B _3505_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_524 VGND VPWR sky130_fd_sc_hd__fill_2
X_2513_ _2159_/A _2513_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3493_ _3504_/A _3491_/Y _3493_/C _4424_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA_clkbuf_4_5_0_clk_i_A clkbuf_4_5_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2444_ _2443_/A _2444_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3226__C _3225_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_229 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2697__C1 _2696_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2375_ _2379_/A _2375_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_644 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3523__A _3514_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_305 VGND VPWR sky130_fd_sc_hd__fill_1
X_4114_ _3974_/A _4039_/B _4033_/A _4113_/X _4576_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_29_519 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_485 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_541 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_530 VGND VPWR sky130_fd_sc_hd__decap_4
X_4045_ _4030_/X _4073_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_83_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_511 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4430__CLK _4430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_393 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_219 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_268 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4504__D _4504_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4073__B _4071_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4580__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_290 VGND VPWR sky130_fd_sc_hd__decap_12
X_3829_ utmi_rxvalid_i _3822_/Y utmi_rxactive_i _3829_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_20_463 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3716__A2 _4474_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2602__A _2601_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3417__B _2763_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_590 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_110 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3433__A _3462_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2991__B _2991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_680 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4264__A _3399_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_213 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4504__RESET_B _2290_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3404__A1 _4240_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4414__D _4414_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_88 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__A outport_data_o[5] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2512__A _2159_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_549 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_684 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_463 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4453__CLK _4450_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_113 VGND VPWR sky130_fd_sc_hd__decap_8
X_2160_ _2163_/A _2160_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4158__B _4153_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_647 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3997__B _3994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4174__A _4188_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_2993_ _2920_/B _2992_/Y _2993_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_61_374 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4324__D _4324_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3946__A2 _3944_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3518__A _2864_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3614_ outport_data_o[7] _3587_/X _3615_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2422__A _2419_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4594_ _4204_/X _4281_/A _2183_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3545_ _3545_/A _3543_/Y _3545_/C _3545_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_115_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_3476_ _3506_/A _3479_/B _3477_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_103_538 VGND VPWR sky130_fd_sc_hd__decap_8
X_2427_ _2431_/A _2427_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4123__A2 _4122_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3253__A _3253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3882__A1 _4539_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2358_ _2358_/A _2358_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_28_38 VGND VPWR sky130_fd_sc_hd__decap_4
X_2289_ _2288_/X _2289_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_5_9_0_clk_i_A clkbuf_5_9_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_617 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_179 VGND VPWR sky130_fd_sc_hd__fill_2
X_4028_ _4562_/Q _4027_/X _4031_/B VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_71_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_15 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4084__A utmi_data_out_o[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_374 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_205 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_569 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_558 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_65 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3428__A _3498_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4326__CLK _4423_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_282 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2332__A _2337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_415 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_74 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4476__CLK _4473_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2986__B _2986_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4114__A2 _4039_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_621 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4259__A _4236_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3322__B1 _2905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_676 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4409__D _4409_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_455 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_658 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_99 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_500 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3610__B _3610_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_661 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2507__A _2504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_544 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_514 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_536 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3389__B1 _3367_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_70 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_569 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_608 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_7 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2242__A _2241_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_297 VGND VPWR sky130_fd_sc_hd__decap_4
X_3330_ _3327_/Y _2860_/C _3329_/X _3330_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_112_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2896__B _4375_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3261_ _3265_/A _3261_/B _3261_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4169__A _4188_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3073__A _3110_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3504__C _3504_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3864__A1 _4531_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_2212_ _2210_/X _2212_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3192_ _2999_/X _3191_/X _3193_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_66_444 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4319__D _2837_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3801__A _3707_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_617 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4497__RESET_B _2299_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3520__B _3518_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_296 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4426__RESET_B _2384_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_371 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3077__C1 _3076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2417__A _2396_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_683 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_171 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4574__SET_B _2206_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_536 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4349__CLK _4325_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2976_ _3289_/A _2972_/A _2975_/Y _2976_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_108_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3248__A _3248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2152__A _2252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_630 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4499__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_4577_ _4134_/Y _2555_/A _2203_/X _4596_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_1_407 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_3528_ _3528_/A _3528_/B _3528_/C _3528_/D _3544_/B VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_89_547 VGND VPWR sky130_fd_sc_hd__fill_2
X_3459_ _3660_/A _3483_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_569 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4079__A _4079_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_219 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3304__B1 _3302_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_591 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3711__A _3713_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_25 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2327__A _2330_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_31 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2815__C1 _2814_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4245__C _4245_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_650 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_480 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_694 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_683 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4208__A2_N _2721_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4032__A1 _4010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4261__B _4261_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3158__A _3154_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2997__A _2849_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_633 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2897__A2 _2880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3605__B _3603_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_87 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_539 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3846__A1 _2645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_433 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3621__A _3617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_617 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4590__RESET_B _2187_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3340__B _3329_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_499 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_691 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2237__A _2236_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_244 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_469 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_683 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4155__C _4154_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_363 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_480 VGND VPWR sky130_fd_sc_hd__decap_8
X_2830_ _2846_/B inport_accept_o VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3994__C _4557_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_322 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4023__B2 _3976_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2761_ _2761_/A _2731_/X _2761_/C _2760_/X _2761_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__4171__B _4169_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3068__A _3067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_416 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_405 VGND VPWR sky130_fd_sc_hd__fill_1
X_2692_ _2620_/B _2810_/B _2692_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4500_ _4500_/D _4500_/Q _2294_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_61_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4602__D _4602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_562 VGND VPWR sky130_fd_sc_hd__fill_2
X_4431_ _3458_/Y _3455_/A _2377_/X _4430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_6_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_600 VGND VPWR sky130_fd_sc_hd__fill_2
X_4362_ _3390_/Y _3388_/A _2459_/X _4388_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3515__B _3512_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_709 VGND VPWR sky130_fd_sc_hd__fill_2
X_3313_ _3317_/A _3312_/Y _3313_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4293_ _4616_/Q _3657_/D _4247_/A _4293_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_112_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_208 VGND VPWR sky130_fd_sc_hd__decap_6
X_3244_ _2849_/A _3244_/B _3251_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4607__RESET_B _2168_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3531__A _3544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_477 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_466 VGND VPWR sky130_fd_sc_hd__decap_4
X_3175_ _3153_/D _3165_/X _3167_/X _3175_/D _3181_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_27_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_105 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_639 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3250__B _3249_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_683 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_672 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_28 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4014__B2 _4066_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2959_ _4328_/Q _2918_/B _2958_/Y _3257_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3773__B1 _3720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4512__D _4513_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_17_0_clk_i_A clkbuf_4_8_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3128__D _3128_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_600 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2610__A _2610_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_208 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3144__C _3381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3828__B2 _3827_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_720 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4348__RESET_B _2477_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4514__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3441__A _3506_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_583 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4256__B _4263_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_244 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3160__B _3141_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3056__A2 _3026_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_300 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_16_0_clk_i clkbuf_4_8_0_clk_i/X _4323_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_41_642 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4272__A _4234_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_355 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clk_i_A clkbuf_2_1_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4422__D _4422_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3764__B1 _3669_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3616__A _3426_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_471 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2520__A _4446_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_576 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_614 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_517 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3054__C _3011_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3819__A1 _2650_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_561 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3295__A2 _3293_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_230 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_436 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4166__B _4163_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4244__B2 _3399_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_661 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_182 VGND VPWR sky130_fd_sc_hd__fill_2
X_3931_ _3931_/A _4041_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_3862_ _4530_/Q _3855_/X _3861_/X _4530_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__4182__A _4182_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_141 VGND VPWR sky130_fd_sc_hd__fill_2
X_2813_ _2694_/A _2633_/X _2810_/B _2813_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_31_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3755__B1 _3719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4332__D _4332_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3793_ _2522_/X _3782_/X _3790_/X _4527_/Q _3792_/X _4486_/D VGND VPWR sky130_fd_sc_hd__a32o_4
X_2744_ _4468_/Q _4219_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__3526__A _3514_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2675_ _2645_/X _2649_/Y _2675_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4414_ _4414_/D _4414_/Q _2398_/X _4410_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__2430__A _2431_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_642 VGND VPWR sky130_fd_sc_hd__fill_2
X_4345_ _4345_/D _3182_/A _2480_/X _4325_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__4537__CLK _4545_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_517 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_102 VGND VPWR sky130_fd_sc_hd__decap_4
X_4276_ _2516_/X _4276_/B _4275_/Y _4614_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__4441__RESET_B _2365_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3261__A _3265_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_241 VGND VPWR sky130_fd_sc_hd__decap_3
X_3227_ _3381_/A _3375_/A _3011_/X _3227_/D _3227_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_82_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_285 VGND VPWR sky130_fd_sc_hd__fill_2
X_3158_ _3154_/X _3158_/B _3156_/X _3158_/D _3158_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_27_414 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4507__D _2683_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_575 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4235__B2 _4257_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3089_ _3043_/X _3088_/Y _3055_/X _3089_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_42_439 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2797__A1 _2788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_130 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2605__A _2604_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3746__B1 _3739_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2549__A1 _2519_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2549__B2 _2548_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3436__A _3431_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2978__C _2974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2340__A _2345_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4529__RESET_B _2261_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_452 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_163 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4267__A _4267_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3171__A _3171_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3602__C _3601_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4417__D _3526_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_406 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4226__B2 _4207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2515__A _2628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_653 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3985__B1 _3921_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3049__C _4354_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2250__A _2248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2960__B2 _3257_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2460_ _2425_/A _2460_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_3_5_0_clk_i_A clkbuf_2_2_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_290 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4478__SET_B _2321_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3065__B _3369_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2391_ _2391_/A _2391_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_303 VGND VPWR sky130_fd_sc_hd__decap_12
X_4130_ _4316_/Q _3960_/B _4231_/C _4130_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_96_634 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_111 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_550 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4177__A _4186_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4061_ _4061_/A _4059_/X _4061_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3081__A _3055_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_199 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_211 VGND VPWR sky130_fd_sc_hd__decap_3
X_3012_ _3007_/X _3008_/X _3010_/X _3011_/X _3012_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__4327__D _4327_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_380 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_266 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4217__A1 _4214_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_480 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2425__A _2425_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3914_ _2571_/X _3913_/Y _2571_/X _4569_/Q _3914_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__3728__B1 _3674_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3845_ _4531_/Q _3844_/X _3845_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_667 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_3776_ _3681_/X _3771_/X _3681_/X _3771_/X _3776_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_2727_ outport_accept_i _2725_/Y _3657_/D _2727_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_9_690 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3256__A _3268_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2160__A _2163_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_238 VGND VPWR sky130_fd_sc_hd__fill_2
X_2658_ _4525_/Q _2658_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_87_601 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_2589_ _2579_/X _2572_/X _2582_/X _2588_/Y _2589_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_4328_ _4328_/D _4328_/Q _2500_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_293 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_455 VGND VPWR sky130_fd_sc_hd__fill_2
X_4259_ _4236_/Y _4263_/B _4261_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_59_358 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_347 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3259__A2 _3257_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3422__C _3422_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_200 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_542 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_372 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3141__D _3128_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4102__A1_N _3915_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4208__B2 _4207_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_36 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_556 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2335__A _2337_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3967__B1 _2552_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_450 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_601 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_483 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_133 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_500 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2989__B _2986_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_126 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3195__A1 _3366_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_599 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4363__RESET_B _2458_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_354 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_398 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_604 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3613__B _3610_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_626 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_114 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3332__C _3332_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_380 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_520 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_309 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_575 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12_0_clk_i_A clkbuf_3_6_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_225 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2245__A _2238_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3326__A1_N _3347_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3958__B1 _2552_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_80 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4163__C _4163_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4080__C1 _4079_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3973__A3 _3971_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3630_ _3415_/Y _3662_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4382__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3561_ _3503_/A _3582_/B _3561_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4610__D _4265_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VPWR sky130_fd_sc_hd__decap_6
X_2512_ _2159_/A _2512_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_671 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_660 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3507__C _3507_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_547 VGND VPWR sky130_fd_sc_hd__fill_2
X_3492_ _3522_/A _3486_/B _3493_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_6_682 VGND VPWR sky130_fd_sc_hd__fill_2
X_2443_ _2443_/A _2443_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3804__A _2601_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2697__B1 _2694_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2374_ _2339_/A _2379_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3523__B _3521_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9_0_clk_i_A clkbuf_4_9_0_clk_i/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4113_ _4109_/X _4111_/X _4112_/Y _4113_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_56_328 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_4044_ _4022_/X _4037_/X _4033_/X _4043_/Y _4564_/D VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_37_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_704 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_586 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_556 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2155__A _2155_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4073__C _4072_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3828_ _3822_/Y _3827_/X _4514_/Q _3827_/X _3828_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_503 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4520__D _3838_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3759_ _3759_/A _3770_/B _3759_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3417__C _2763_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_517 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_464 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_263 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_497 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_615 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_520 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_531 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_607 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_523 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4264__B _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_578 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3404__A2 _3386_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_67 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4280__A _2516_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4544__RESET_B _2242_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_330 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__B _3592_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_43 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4430__D _3454_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_652 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4117__B1 _3987_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3624__A _4379_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_7 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_475 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_434 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_467 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_564 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3997__C _4558_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4605__D _4605_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4174__B _4169_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2992_ _2944_/Y _2985_/X _2988_/Y _2991_/X _2992_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_34_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2603__B1 _2602_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_291 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3946__A3 _3945_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_127 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4190__A _4620_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2703__A _2702_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3518__B _3512_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3613_ _4393_/Q _3610_/B _3613_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4340__D _3313_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4593_ _4593_/D _4620_/D _2184_/X _4595_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3544_ _3516_/A _3544_/B _3545_/C VGND VPWR sky130_fd_sc_hd__and2_4
X_3475_ _2900_/A _3478_/B _3475_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_103_506 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3534__A _4403_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_2426_ _2431_/A _2426_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3253__B _2956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3882__A2 _3869_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_464 VGND VPWR sky130_fd_sc_hd__fill_2
X_2357_ _2358_/A _2357_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_306 VGND VPWR sky130_fd_sc_hd__decap_4
X_2288_ _2253_/A _2288_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_309 VGND VPWR sky130_fd_sc_hd__decap_6
X_4027_ _3957_/Y _4026_/X _3957_/Y _4026_/X _4027_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_372 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_512 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4515__D _3829_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4084__B _4082_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_556 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4044__C1 _4043_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_548 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3709__A _3713_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_15 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3428__B _3428_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_182 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_377 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3444__A outport_data_o[2] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4259__B _4263_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3322__A1 _2849_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_644 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_572 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3322__B2 _3321_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3694__A2_N _3693_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_78 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_489 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_478 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_61 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_383 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4425__D _4425_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_342 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2833__B1 _2832_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_567 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_386 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4035__C1 _4034_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3389__A1 _3388_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_60 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3619__A _3640_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2523__A _4487_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_93 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_119 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4420__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_504 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_314 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2896__C _2895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3354__A _3353_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_460 VGND VPWR sky130_fd_sc_hd__fill_2
X_3260_ _3268_/A _3260_/B _4328_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_3_493 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_482 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4169__B _4167_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_412 VGND VPWR sky130_fd_sc_hd__decap_12
X_3191_ _3136_/X _3176_/X _3191_/C _3190_/X _3191_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_2211_ _2210_/X _2211_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3864__A2 _3855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_659 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4570__CLK _4323_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3801__B _2639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4185__A _4185_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_350 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3520__C _3520_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_275 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_415 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3077__B1 _3074_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2824__B1 _2796_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4335__D _3292_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4466__RESET_B _2335_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_548 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3529__A _3544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2433__A _2434_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2975_ _2933_/X _2975_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_30_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3772__A1_N _3695_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3001__B1 _2850_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4576_ _4576_/D _3974_/A _2204_/X _4574_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_116_642 VGND VPWR sky130_fd_sc_hd__decap_4
X_3527_ _3508_/A _3545_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3264__A _3268_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_526 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_358 VGND VPWR sky130_fd_sc_hd__fill_2
X_3458_ _3424_/X _3458_/B _3457_/X _3458_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3304__A1 _3280_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_38 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4079__B _4079_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2409_ _2408_/A _2409_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_570 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3304__B2 _3248_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3389_ _3388_/Y _3386_/X _3367_/A _3389_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_69_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_423 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3711__B _3711_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_37 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2608__A _2566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_448 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2815__B1 _2811_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_43 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4245__D _4244_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_515 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_397 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3439__A _4427_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1_0_clk_i_A clkbuf_0_clk_i/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_356 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4032__A2 _4031_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2343__A _2345_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2981__A1_N _4429_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4261__C _4261_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3158__B _3158_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4443__CLK _4446_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_664 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2997__B _2915_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_11 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_12_0_clk_i clkbuf_4_6_0_clk_i/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__3174__A _3220_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4593__CLK _4595_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_645 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3605__C _3604_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_507 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3902__A utmi_data_in_i[4] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3846__A2 _3841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_437 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_70 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_673 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3349__A _3397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2253__A _2253_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2760_ _4497_/Q _2730_/X _2760_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4171__C _4170_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_581 VGND VPWR sky130_fd_sc_hd__fill_2
X_2691_ _2691_/A _2691_/B _2691_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_428 VGND VPWR sky130_fd_sc_hd__fill_2
X_4430_ _3454_/Y _3451_/A _2378_/X _4430_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_8_596 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_64 VGND VPWR sky130_fd_sc_hd__decap_4
X_4361_ _4361_/D _4361_/Q _2461_/X _4334_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3084__A _3084_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_122 VGND VPWR sky130_fd_sc_hd__fill_1
X_3312_ _3251_/A _3310_/X _3311_/X _2986_/A _3248_/A _3312_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_4292_ _4283_/Y _4284_/X _4291_/Y _4292_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_113_689 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_177 VGND VPWR sky130_fd_sc_hd__decap_12
X_3243_ _2954_/Y _3243_/B _3243_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_66_220 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3812__A _3812_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_242 VGND VPWR sky130_fd_sc_hd__decap_12
X_3174_ _3220_/C _3174_/B _3171_/X _3173_/X _3175_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_82_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2428__A _2431_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_286 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_489 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4316__CLK _4612_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_459 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4466__CLK _4497_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2958_ _2920_/B _2958_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2163__A _2163_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_389 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3773__A1 _3769_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2889_ _3367_/A _2996_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_612 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_216 VGND VPWR sky130_fd_sc_hd__decap_12
X_4559_ _4001_/Y _4559_/Q _2225_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_103_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_356 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3144__D _3008_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3722__A _3670_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_76 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3441__B _3437_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4388__RESET_B _2429_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_426 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2338__A _2381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_448 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3160__C _3216_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_289 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_256 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4317__RESET_B _2512_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_662 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_68 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4272__B _4253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_665 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3213__B1 _3212_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_327 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3764__B2 _3763_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2801__A _2801_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3616__B _3427_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_529 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3054__D _3010_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_497 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_626 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3819__A2 _3804_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3632__A outport_data_o[3] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4339__CLK _4430_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_710 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3295__A3 _3294_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2248__A _2248_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4489__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_576 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_418 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_651 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_109 VGND VPWR sky130_fd_sc_hd__decap_12
X_3930_ _2604_/X _3927_/Y _3928_/X _2581_/A _3929_/Y _3930_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_32_632 VGND VPWR sky130_fd_sc_hd__fill_2
X_3861_ _4538_/Q _3859_/B _3861_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__3079__A _3350_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_654 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_665 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_676 VGND VPWR sky130_fd_sc_hd__fill_2
X_3792_ _3792_/A _3792_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_82_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_2812_ _2796_/B _2799_/A _2812_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__4613__D _4274_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_715 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3755__A1 _3726_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2743_ _2743_/A _4443_/Q _2743_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_117_258 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_2674_ _4524_/Q _2674_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2711__A _2710_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4413_ _3514_/Y _4413_/Q _2399_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3526__B _3524_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_420 VGND VPWR sky130_fd_sc_hd__decap_3
X_4344_ _4344_/D _3161_/A _2481_/X _4325_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_453 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_615 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_604 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_676 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_142 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3542__A _3545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_348 VGND VPWR sky130_fd_sc_hd__fill_2
X_4275_ _4497_/Q _2761_/A _3657_/D _4213_/Y _4614_/Q _4275_/Y VGND VPWR sky130_fd_sc_hd__a41oi_4
XANTENNA__3261__B _3261_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_136 VGND VPWR sky130_fd_sc_hd__fill_2
X_3226_ _3397_/A _3216_/X _3225_/Y _3226_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_82_510 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2158__A _2252_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3157_ _3059_/Y _3094_/X _3055_/X _3158_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_94_381 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_437 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4410__RESET_B _2402_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_109 VGND VPWR sky130_fd_sc_hd__decap_12
X_3088_ _3087_/X _3088_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_35_470 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2797__A2 _2796_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4523__D _3846_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3746__B2 _3745_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_704 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3746__A1 _3671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_495 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2549__A2 _2547_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_348 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3717__A _3717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_247 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2621__A _2601_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2978__D _2978_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3452__A outport_data_o[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4267__B _4264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_318 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_595 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_724 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3171__B _3171_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3131__C1 _2997_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3682__B1 _3668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_705 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4283__A _2533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_632 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3985__A1 _3984_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3985__B2 _3981_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4433__D _3467_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_153 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_164 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_157 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3627__A _2880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3049__D _3120_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2531__A _2524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_385 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3065__C _3046_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2390_ _2391_/A _2390_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_122_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_646 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_315 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3362__A _3397_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_348 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_540 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4177__B _4178_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_98 VGND VPWR sky130_fd_sc_hd__fill_2
X_4060_ _4061_/A _4059_/X _4062_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_95_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_90 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4608__D _4608_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_573 VGND VPWR sky130_fd_sc_hd__fill_2
X_3011_ _4358_/Q _3011_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3081__B _3080_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_532 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4217__A2 _4216_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_226 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2706__A _2706_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4193__A _4197_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3913_ _2604_/X _3910_/Y _3911_/X _2581_/A _3912_/Y _3913_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_3844_ _3824_/X _3844_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4343__D _3133_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_646 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3537__A _4404_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3728__B2 _3727_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3775_ _3724_/A _3673_/A _2687_/X _3774_/X _3775_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_118_556 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2441__A _2443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4504__CLK _4486_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_2726_ _3417_/D _3657_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_578 VGND VPWR sky130_fd_sc_hd__fill_2
X_2657_ _4521_/Q _2657_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3256__B _3256_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_451 VGND VPWR sky130_fd_sc_hd__fill_2
X_2588_ _2581_/X _2587_/Y _2588_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3272__A _3268_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_473 VGND VPWR sky130_fd_sc_hd__fill_2
X_4327_ _4327_/D _2917_/A _2501_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_86_101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_315 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_657 VGND VPWR sky130_fd_sc_hd__fill_2
X_4258_ _4265_/A _4258_/B _4258_/C _4608_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_47_27 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4518__D _4518_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3259__A3 _3258_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_489 VGND VPWR sky130_fd_sc_hd__fill_2
X_3209_ _3209_/A _3205_/X _3208_/X _3179_/Y _3209_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_103_33 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3664__B1 _3663_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4189_ _4182_/Y _4186_/X _4187_/X _4189_/D _4202_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_55_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_48 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3967__A1 _2579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3967__B2 _3966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4484__SET_B _2314_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3447__A _4429_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2351__A _2352_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3195__A2 _2916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_602 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4278__A _2537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_388 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3182__A _3182_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_123 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4332__RESET_B _2495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4428__D _3446_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3332__D _2872_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_329 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3910__A _4317_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_159 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_565 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_82 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2526__A _2522_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_579 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3958__B2 _3957_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3958__A1 _2578_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4080__B1 _4050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4527__CLK _4534_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_270 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2261__A _2261_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3560_ _3583_/B _3582_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_2511_ _2159_/A _2511_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_559 VGND VPWR sky130_fd_sc_hd__fill_2
X_3491_ _3491_/A _3479_/B _3491_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_5_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_2442_ _2443_/A _2442_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_602 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_193 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3894__B1 _3893_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_421 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2697__A1 _2687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3804__B _3804_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_635 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4188__A _4153_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2373_ _2367_/X _2373_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3092__A _3176_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3523__C _3523_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_145 VGND VPWR sky130_fd_sc_hd__decap_8
X_4112_ _4109_/X _4111_/X _4030_/X _4112_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_110_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_178 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_167 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4338__D _3305_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4043_ _4043_/A _4039_/B _4043_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3820__A _3820_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_19 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_660 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2436__A _2434_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_524 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_281 VGND VPWR sky130_fd_sc_hd__fill_2
X_3827_ _3883_/A _3827_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4070__A2_N _4069_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_342 VGND VPWR sky130_fd_sc_hd__fill_2
X_3758_ _3759_/A _3770_/B _3760_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__2171__A _2168_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2709_ _4499_/Q _3806_/A _4502_/Q _3816_/A _2730_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_4_609 VGND VPWR sky130_fd_sc_hd__fill_2
X_3689_ _4520_/Q _2657_/X _2643_/Y _2641_/Y _3691_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__3417__D _3417_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4126__A1 _4123_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_581 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3885__B1 _3884_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_476 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3730__A _3730_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_649 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_87 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_619 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_502 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2346__A _2339_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4023__A2_N utmi_data_out_o[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_226 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_557 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_719 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_590 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4280__B _4276_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_454 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_465 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3177__A _3110_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_33 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4584__RESET_B _2194_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4117__A1 _3987_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4513__RESET_B _2279_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_207 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4117__B2 _3999_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_570 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_229 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3624__B _3620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3876__B1 _3875_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_454 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3640__A _4384_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_619 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2256__A _2258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_535 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_513 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_598 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_395 VGND VPWR sky130_fd_sc_hd__fill_2
X_2991_ _3464_/A _2991_/B _2991_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_61_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3800__B1 _2659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2603__A1 _3993_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_75 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4190__B _4202_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_3612_ _3612_/A _3610_/X _3611_/X _4392_/D VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__3087__A _3086_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4592_ _4592_/D _4592_/Q _2185_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3543_ _3543_/A _3543_/B _3543_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_367 VGND VPWR sky130_fd_sc_hd__fill_2
X_3474_ _3483_/A _3471_/Y _3473_/X _3474_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_89_708 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_491 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3534__B _3543_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_529 VGND VPWR sky130_fd_sc_hd__decap_6
X_2425_ _2425_/A _2431_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_432 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_421 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_573 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_240 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_402 VGND VPWR sky130_fd_sc_hd__decap_3
X_2356_ _2358_/A _2356_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_28_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_595 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3550__A _2865_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_435 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_424 VGND VPWR sky130_fd_sc_hd__fill_2
X_2287_ _2283_/A _2287_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_660 VGND VPWR sky130_fd_sc_hd__decap_8
X_4026_ _4099_/B _4025_/X _4099_/B _4025_/X _4026_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4292__B1 _4291_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2166__A _2252_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_652 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_181 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_568 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4044__B1 _4033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3709__B _3709_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4531__D _3864_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_651 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_43 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_326 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3322__A2 _3319_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_562 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_627 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_595 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4372__CLK _4551_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3460__A _3460_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_438 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_129 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_107 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_671 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_170 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_449 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2833__A1 _4317_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_685 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4035__B1 _4033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_527 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2804__A _2804_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_195 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3389__A2 _3386_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_83 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_240 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_284 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4441__D _2723_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_266 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_161 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3635__A outport_data_o[4] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3354__B _2857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_2210_ _2238_/A _2210_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_3190_ _3074_/X _3189_/Y _3190_/C _3165_/X _3190_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_120_381 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_370 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_210 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_424 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3077__A1 _3059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_438 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4616__D _4616_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2824__B2 _2823_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2824__A1 _2821_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_343 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_395 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4026__B1 _4099_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2974_ _2902_/D _2973_/X _2902_/D _2973_/X _2974_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_61_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2714__A _2587_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_590 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4351__D _3004_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_560 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4435__RESET_B _2372_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_593 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3001__A1 _2886_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4575_ _4107_/X _3964_/A _2205_/X _4574_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA__3545__A _3545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_142 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_3526_ _3514_/A _3524_/Y _3525_/X _3526_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_89_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_698 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3264__B _3264_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_197 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4395__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_3457_ _3547_/A _3462_/B _3457_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_39_28 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4079__C _4079_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_2408_ _2408_/A _2408_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3304__A2 _3302_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3388_ _3388_/A _3388_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_2339_ _2339_/A _2345_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3280__A _3251_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_446 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_608 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4526__D _3852_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_107 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2608__B _2607_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4009_ _3933_/Y _4565_/Q _4563_/Q _3949_/Y _4009_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_111_22 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2815__A1 _2788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_66 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2624__A _2624_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_527 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3439__B _3434_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2963__A2_N _3261_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3158__C _3156_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4008__A1_N _4569_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_120 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3455__A _3455_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_602 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3174__B _3174_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_63 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_464 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3902__B _3904_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4286__A _3808_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_413 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_497 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3190__A _3074_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4436__D _4436_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4008__B1 _4569_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2534__A _2533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_398 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3349__B _3345_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_7 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3231__A1 _2916_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_520 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2690_ _3707_/A _3720_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_4360_ _4360_/D _4360_/Q _2462_/X _4334_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_98_313 VGND VPWR sky130_fd_sc_hd__fill_2
X_3311_ _3253_/A _2987_/X _3311_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2742__B1 _2736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_657 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_646 VGND VPWR sky130_fd_sc_hd__fill_1
X_4291_ _2548_/A _2761_/A _2533_/X _4288_/Y _4290_/X _4291_/Y VGND VPWR sky130_fd_sc_hd__o32ai_4
XFILLER_112_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_368 VGND VPWR sky130_fd_sc_hd__fill_1
X_3242_ _3265_/A _3243_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_402 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_189 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_593 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3812__B _3805_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2709__A _4499_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3173_ _3041_/X _3172_/X _3095_/X _3122_/Y _3173_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__4196__A _4194_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_232 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_574 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_416 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_619 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4346__D _3193_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_298 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_663 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_652 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2444__A _2443_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_493 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_622 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_696 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4616__RESET_B _2155_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_346 VGND VPWR sky130_fd_sc_hd__fill_2
X_2957_ _2900_/A _2956_/X _2900_/A _2956_/X _2957_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_41_29 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_18 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3773__A2 _3772_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2888_ _3392_/A _3367_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3693__A2_N _3692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2981__B1 _4429_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3275__A _2926_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4558_ _4558_/D _4558_/Q _2226_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3509_ _4412_/Q _3512_/B _3509_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_103_123 VGND VPWR sky130_fd_sc_hd__fill_2
X_4489_ _4489_/D _4489_/Q _2308_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_1_228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_519 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_690 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3722__B _3723_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_541 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2619__A _2618_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_202 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4238__B1 _4237_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3160__D _3160_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_674 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4410__CLK _4410_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_58 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2354__A _2358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_110 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4357__RESET_B _2465_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_52 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_154 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3213__A1 _2999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_339 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4560__CLK _4560_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_523 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_51 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_534 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3185__A _4346_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3616__C _3528_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_495 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_508 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_638 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3632__B _3625_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_722 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_530 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_416 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_588 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_3860_ _4529_/Q _3855_/X _3859_/X _4529_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__2264__A _2261_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3156__A1_N _3029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_121 VGND VPWR sky130_fd_sc_hd__fill_1
X_3791_ _3785_/A _3792_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2811_ _2699_/X _2810_/X _3704_/A _2811_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__3079__B _4357_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3755__A2 _3713_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VPWR sky130_fd_sc_hd__decap_8
X_2742_ _2738_/X _2741_/X _2736_/X _2742_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_12_390 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2963__B1 _4421_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_4412_ _4412_/D _4412_/Q _2400_/X _4331_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2673_ _4520_/Q _2673_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3095__A _3048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_383 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3526__C _3525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_611 VGND VPWR sky130_fd_sc_hd__fill_2
X_4343_ _3133_/Y _3005_/A _2483_/X _4325_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3823__A utmi_rxactive_i VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_443 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_165 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_4274_ _2516_/X _4272_/X _4273_/Y _4274_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__3542__B _3542_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_498 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_476 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_638 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_627 VGND VPWR sky130_fd_sc_hd__decap_4
X_3225_ _3077_/X _3221_/X _3224_/X _3202_/C _3225_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_67_541 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_530 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2439__A _2425_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4433__CLK _4418_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_574 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_265 VGND VPWR sky130_fd_sc_hd__decap_4
X_3156_ _3029_/X _3070_/X _3066_/A _3036_/X _3156_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_3087_ _3086_/X _3087_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_82_555 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_599 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_482 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_633 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4450__RESET_B _2355_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4583__CLK _4596_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2174__A _2166_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_644 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_474 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3746__A2 _4474_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2902__A _3488_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3989_ _2701_/A _3988_/X _4555_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_108_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3717__B _3674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_548 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_487 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_349 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2349__A _2352_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_541 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3131__B1 _3130_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_585 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_563 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3171__C _3130_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3682__B2 _3675_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_393 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_522 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_235 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4538__RESET_B _2249_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_419 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_227 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4283__B _4283_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_622 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_84 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3985__A2 _3979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_463 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_688 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3908__A utmi_data_in_i[7] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2812__A _2796_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_50 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3198__B1 _3085_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3627__B _3620_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_708 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2531__B _2531_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_397 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_375 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3065__D _3375_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3643__A _3643_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3370__B1 _3369_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_273 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_424 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_327 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4456__CLK _4509_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3362__B _3358_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_457 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2259__A _2258_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_468 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_500 VGND VPWR sky130_fd_sc_hd__fill_2
X_3010_ _3009_/Y _3010_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_91_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_544 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_385 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_205 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2706__B _2910_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4193__B _4196_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3912_ _4553_/Q _3912_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3843_ _3685_/X _3841_/X _3842_/X _3843_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_32_463 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3818__A _3818_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2722__A _2721_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3537__B _3543_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_3774_ _3769_/X _3772_/X _3773_/Y _3774_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_2725_ _4489_/Q _4488_/Q _2527_/Y _2525_/X _2725_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
X_2656_ _2696_/A _2633_/X _2655_/X _2671_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__3553__A _2865_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2587_ _4316_/Q _3960_/B _4342_/Q _3417_/D _2587_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XANTENNA__3272__B _3271_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4326_ _3250_/Y _2917_/B _2502_/X _4423_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_87_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_4257_ _4257_/A _4264_/B _4258_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__2169__A _2168_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4188_ _4153_/A _4153_/B _4188_/C _4188_/D _4189_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_3208_ _3208_/A _3176_/X _3206_/X _3207_/X _3208_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_28_703 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3664__A1 _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_382 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_533 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_522 VGND VPWR sky130_fd_sc_hd__fill_2
X_3139_ _3059_/Y _3150_/D _3188_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_55_577 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_566 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_419 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4534__D _3871_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3967__A2 _3965_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_260 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4329__CLK _4331_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_124 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_636 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_658 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2632__A _2784_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3447__B _3434_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_97 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4479__CLK _4470_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3463__A _3483_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4278__B _2730_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_284 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_703 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_714 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_691 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3910__B _2585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4372__RESET_B _2448_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2807__A _2691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_94 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_717 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_374 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2526__B _2525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_547 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4444__D _2742_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3958__A2 _3956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4080__A1 _3931_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_452 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3638__A outport_data_o[5] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2542__A _4498_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_3490_ _3504_/A _3488_/Y _3490_/C _4423_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_2510_ _2159_/A _2510_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_2441_ _2443_/A _2441_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3343__B1 _3332_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_722 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3894__A1 _4544_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2697__A2 _2689_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4188__B _4153_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2372_ _2367_/X _2372_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_135 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4619__D _4619_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_4111_ _4026_/X _4110_/X _4026_/X _4110_/X _4111_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__3092__B _3059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_254 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_308 VGND VPWR sky130_fd_sc_hd__decap_3
X_4042_ _4563_/Q _4037_/X _4033_/X _4041_/Y _4042_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_110_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3820__B _3804_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_522 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2717__A _2761_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_374 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4354__D _3339_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_290 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3548__A _3545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_433 VGND VPWR sky130_fd_sc_hd__decap_4
X_3826_ _3904_/B _3883_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__2452__A _2449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_332 VGND VPWR sky130_fd_sc_hd__decap_4
X_3757_ _3683_/A _3668_/X _3667_/A _3668_/A _3770_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_2708_ _4503_/Q _3816_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_387 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_376 VGND VPWR sky130_fd_sc_hd__fill_2
X_3688_ _4524_/Q _4525_/Q _2674_/Y _2658_/Y _3690_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_3_109 VGND VPWR sky130_fd_sc_hd__fill_2
X_2639_ _2638_/Y _2639_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4126__A2 _4125_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3885__A1 _4540_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4529__D _4529_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_221 VGND VPWR sky130_fd_sc_hd__fill_2
X_4309_ _2159_/A _4309_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_606 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3730__B _3730_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_511 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2627__A _2626_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_514 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_588 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_599 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_388 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_208 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3458__A _3424_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4280__C _4280_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2362__A _2362_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_415 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_444 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_41 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_477 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3177__B _3363_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_56 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4117__A2 _4602_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3193__A _2996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3876__A1 _4536_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_665 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4439__D _4439_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_414 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_105 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4553__RESET_B _2232_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3921__A _4554_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_425 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3640__B _3640_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4563__SET_B _2220_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2537__A _4500_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_81 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2764__A1_N _4234_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2990_ _3314_/A _2986_/Y _2989_/X _2991_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_9_10 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3800__A1 _2601_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3800__B2 _3792_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2603__A2 _2599_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2272__A _2272_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3611_ outport_data_o[6] _3587_/X _3611_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_80_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_98 VGND VPWR sky130_fd_sc_hd__fill_2
X_4591_ _4197_/X _4591_/Q _2186_/X _4446_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3542_ _3545_/A _3542_/B _3542_/C _3542_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_3473_ _3503_/A _3479_/B _3473_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__4199__A _4198_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_400 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3316__B1 _3314_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_2424_ _2381_/A _2425_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_2355_ _2358_/A _2355_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__4349__D _3226_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3831__A _4517_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_252 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_606 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3550__B _3541_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_2286_ _2283_/A _2286_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_469 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2447__A _2449_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4292__A1 _4283_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4025_ _4022_/X _4024_/B _4024_/Y _4025_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_65_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_525 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_642 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_536 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_355 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4044__A1 _4022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_388 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_720 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2182__A _2183_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3809_ _2641_/Y _3803_/X _3808_/X _3809_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_20_263 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_407 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_162 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_55 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2910__A _2560_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_602 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4517__CLK _4519_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3322__A3 _3320_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_116 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3460__B _3437_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_469 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_458 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_447 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2357__A _2358_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4238__A1_N _4236_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_653 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2833__A2 _2831_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_536 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_377 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_355 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4035__A1 _4561_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_506 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2804__B _3704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_591 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3794__B1 _2673_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3188__A _3188_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_289 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3635__B _3625_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_349 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_327 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3651__A _3522_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_723 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_639 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2267__A _2253_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_80 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_661 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_672 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3077__A2 _3205_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_491 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2824__A2 _2788_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_642 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4026__B2 _4025_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_2973_ _2930_/A _2948_/A _2972_/Y _2973_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_61_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2714__B _2713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3098__A _3097_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_572 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3826__A _3904_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2730__A _3810_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3001__A2 _2906_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_4574_ _4098_/X _3955_/A _2206_/X _4574_/CLK VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_116_666 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3545__B _3543_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3525_ _3554_/A _3516_/B _3525_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_89_517 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4404__RESET_B _2409_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_338 VGND VPWR sky130_fd_sc_hd__fill_1
X_3456_ outport_data_o[5] _3547_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_2407_ _2408_/A _2407_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_550 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3561__A _3503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3304__A3 _3303_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_3387_ _3386_/X _3394_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_583 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_263 VGND VPWR sky130_fd_sc_hd__fill_2
X_2338_ _2381_/A _2339_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_127 VGND VPWR sky130_fd_sc_hd__decap_4
X_2269_ _2272_/A _2269_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_55_17 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2177__A _2177_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_119 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_160 VGND VPWR sky130_fd_sc_hd__decap_4
X_4008_ _4569_/Q _4007_/X _4569_/Q _4007_/X _4008_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_300 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2815__A2 _2809_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_56 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2905__A _2905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_16 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_539 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3776__B1 _3681_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4542__D _3890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_583 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3736__A _3736_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3158__D _3158_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_482 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_611 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2640__A _2628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_716 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3455__B _3434_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_614 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_699 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_143 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3174__C _3171_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_259 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_86 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3471__A _4418_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_443 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3700__B1 _3682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_712 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4286__B _4498_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_425 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_609 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3190__B _3189_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_247 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_322 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_269 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4008__B2 _4007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_366 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_472 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4100__A1_N _3918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_377 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_9 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4452__D _2681_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3349__C _3349_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_358 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3231__A2 _3228_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_561 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_408 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3646__A _3528_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_71 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2990__A1 _3314_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2550__A _2701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_44 VGND VPWR sky130_fd_sc_hd__decap_3
X_3310_ _2986_/A _3246_/A _3310_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__2742__A1 _2738_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_636 VGND VPWR sky130_fd_sc_hd__fill_2
X_4290_ _2548_/Y _2718_/B _2718_/B _4289_/X _4290_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_113_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_509 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_550 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_701 VGND VPWR sky130_fd_sc_hd__fill_2
X_3241_ _3241_/A _3265_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__3381__A _3381_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_520 VGND VPWR sky130_fd_sc_hd__decap_4
X_3172_ _3110_/C _3018_/X _3172_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4196__B _4196_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_691 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2709__B _3806_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_108 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2725__A _4489_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_483 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_634 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4362__D _3390_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_2956_ _2917_/A _2917_/B _2956_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_22_369 VGND VPWR sky130_fd_sc_hd__fill_2
X_2887_ _2905_/A _2886_/X _2887_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__3556__A _3528_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2981__B2 _3298_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2460__A _2425_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4362__CLK _4388_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_441 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3275__B _3275_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4183__B1 _4182_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_463 VGND VPWR sky130_fd_sc_hd__fill_2
X_4557_ _4557_/D _4557_/Q _2227_/X _4560_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3508_ _3508_/A _3514_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_347 VGND VPWR sky130_fd_sc_hd__fill_2
X_4488_ _3788_/X _4488_/Q _2309_/X _4486_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA__3930__B1 _2581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_669 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_146 VGND VPWR sky130_fd_sc_hd__decap_4
X_3439_ _4427_/Q _3434_/B _3439_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_106_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_380 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4537__D _4537_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_609 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_704 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4238__B2 _4270_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_428 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_620 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2635__A _2635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_656 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_645 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_122 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_336 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_347 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3213__A2 _3209_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4397__RESET_B _2418_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3466__A _3554_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2370__A _2367_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_290 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4326__RESET_B _2502_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_463 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3616__D _3498_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_466 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_273 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4447__D _4447_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_520 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_564 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_523 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_480 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_269 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2545__A _2544_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_664 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3988__B1 _3929_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_2810_ _2636_/A _2810_/B _2810_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3790_ _2669_/A _3790_/B _3790_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__4385__CLK _4380_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3079__C _4354_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_177 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VPWR sky130_fd_sc_hd__decap_3
X_2741_ _2718_/B _2741_/B _2716_/Y _2740_/X _2741_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_12_380 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2963__B2 _3261_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2280__A _2277_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3376__A _3376_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4411_ _3507_/Y _4411_/Q _2401_/X _4410_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_227 VGND VPWR sky130_fd_sc_hd__fill_2
X_2672_ _2785_/C _3780_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_68_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4069__A1_N _3933_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_4342_ _3239_/Y _4342_/Q _2484_/X _4342_/CLK VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_667 VGND VPWR sky130_fd_sc_hd__decap_4
X_4273_ _4368_/Q _4263_/B _4273_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__3542__C _3542_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_317 VGND VPWR sky130_fd_sc_hd__decap_12
X_3224_ _3224_/A _3156_/X _3167_/X _3224_/D _3224_/X VGND VPWR sky130_fd_sc_hd__or4_4
.ends

